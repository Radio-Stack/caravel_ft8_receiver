magic
tech sky130A
magscale 1 2
timestamp 1620311099
<< mvpsubdiff >>
rect 338844 634421 338868 635198
rect 364182 634421 364206 635198
<< mvpsubdiffcont >>
rect 338868 634421 364182 635198
<< locali >>
rect 338852 634421 338868 635198
rect 364182 634421 364198 635198
<< viali >>
rect 350697 634466 352402 635166
<< metal1 >>
rect 350574 635565 352546 635623
rect 350574 634223 350642 635565
rect 352492 634223 352546 635565
rect 350574 634156 352546 634223
<< via1 >>
rect 350642 635166 352492 635565
rect 350642 634466 350697 635166
rect 350697 634466 352402 635166
rect 352402 634466 352492 635166
rect 350642 634223 352492 634466
<< metal2 >>
rect 350574 635565 352546 635623
rect 350574 634223 350642 635565
rect 352492 634223 352546 635565
rect 350574 634156 352546 634223
rect -6372 5366 -6260 6646
rect -5190 5366 -5078 6646
rect -4008 5366 -3896 6646
rect -2826 5366 -2714 6646
rect -1644 5366 -1532 6646
rect -462 5366 -350 6646
rect 720 5366 832 6646
rect 1902 5366 2014 6646
rect 3084 5366 3196 6646
rect 4266 5366 4378 6646
rect 5448 5366 5560 6646
rect 6630 5366 6742 6646
rect 7812 5366 7924 6646
rect 8994 5366 9106 6646
rect 10176 5366 10288 6646
rect 11358 5366 11470 6646
rect 12540 5366 12652 6646
rect 13722 5366 13834 6646
rect 14904 5366 15016 6646
rect 16086 5366 16198 6646
rect 17268 5366 17380 6646
rect 18450 5366 18562 6646
rect 19632 5366 19744 6646
rect 20814 5366 20926 6646
rect 21996 5366 22108 6646
rect 23178 5366 23290 6646
rect 24360 5366 24472 6646
rect 25542 5366 25654 6646
rect 26724 5366 26836 6646
rect 27906 5366 28018 6646
rect 29088 5366 29200 6646
rect 30270 5366 30382 6646
rect 31452 5366 31564 6646
rect 32634 5366 32746 6646
rect 33816 5366 33928 6646
rect 34998 5366 35110 6646
rect 36180 5366 36292 6646
rect 37362 5366 37474 6646
rect 38544 5366 38656 6646
rect 39726 5366 39838 6646
rect 40908 5366 41020 6646
rect 42090 5366 42202 6646
rect 43272 5366 43384 6646
rect 44454 5366 44566 6646
rect 45636 5366 45748 6646
rect 46818 5366 46930 6646
rect 48000 5366 48112 6646
rect 49182 5366 49294 6646
rect 50364 5366 50476 6646
rect 51546 5366 51658 6646
rect 52728 5366 52840 6646
rect 53910 5366 54022 6646
rect 55092 5366 55204 6646
rect 56274 5366 56386 6646
rect 57456 5366 57568 6646
rect 58638 5366 58750 6646
rect 59820 5366 59932 6646
rect 61002 5366 61114 6646
rect 62184 5366 62296 6646
rect 63366 5366 63478 6646
rect 64548 5366 64660 6646
rect 65730 5366 65842 6646
rect 66912 5366 67024 6646
rect 68094 5366 68206 6646
rect 69276 5366 69388 6646
rect 70458 5366 70570 6646
rect 71640 5366 71752 6646
rect 72822 5366 72934 6646
rect 74004 5366 74116 6646
rect 75186 5366 75298 6646
rect 76368 5366 76480 6646
rect 77550 5366 77662 6646
rect 78732 5366 78844 6646
rect 79914 5366 80026 6646
rect 81096 5366 81208 6646
rect 82278 5366 82390 6646
rect 83460 5366 83572 6646
rect 84642 5366 84754 6646
rect 85824 5366 85936 6646
rect 87006 5366 87118 6646
rect 88188 5366 88300 6646
rect 89370 5366 89482 6646
rect 90552 5366 90664 6646
rect 91734 5366 91846 6646
rect 92916 5366 93028 6646
rect 94098 5366 94210 6646
rect 95280 5366 95392 6646
rect 96462 5366 96574 6646
rect 97644 5366 97756 6646
rect 98826 5366 98938 6646
rect 100008 5366 100120 6646
rect 101190 5366 101302 6646
rect 102372 5366 102484 6646
rect 103554 5366 103666 6646
rect 104736 5366 104848 6646
rect 105918 5366 106030 6646
rect 107100 5366 107212 6646
rect 108282 5366 108394 6646
rect 109464 5366 109576 6646
rect 110646 5366 110758 6646
rect 111828 5366 111940 6646
rect 113010 5366 113122 6646
rect 114192 5366 114304 6646
rect 115374 5366 115486 6646
rect 116556 5366 116668 6646
rect 117738 5366 117850 6646
rect 118920 5366 119032 6646
rect 120102 5366 120214 6646
rect 121284 5366 121396 6646
rect 122466 5366 122578 6646
rect 123648 5366 123760 6646
rect 124830 5366 124942 6646
rect 126012 5366 126124 6646
rect 127194 5366 127306 6646
rect 128376 5366 128488 6646
rect 129558 5366 129670 6646
rect 130740 5366 130852 6646
rect 131922 5366 132034 6646
rect 133104 5366 133216 6646
rect 134286 5366 134398 6646
rect 135468 5366 135580 6646
rect 136650 5366 136762 6646
rect 137832 5366 137944 6646
rect 139014 5366 139126 6646
rect 140196 5366 140308 6646
rect 141378 5366 141490 6646
rect 142560 5366 142672 6646
rect 143742 5366 143854 6646
rect 144924 5366 145036 6646
rect 146106 5366 146218 6646
rect 147288 5366 147400 6646
rect 148470 5366 148582 6646
rect 149652 5366 149764 6646
rect 150834 5366 150946 6646
rect 152016 5366 152128 6646
rect 153198 5366 153310 6646
rect 154380 5366 154492 6646
rect 155562 5366 155674 6646
rect 156744 5366 156856 6646
rect 157926 5366 158038 6646
rect 159108 5366 159220 6646
rect 160290 5366 160402 6646
rect 161472 5366 161584 6646
rect 162654 5366 162766 6646
rect 163836 5366 163948 6646
rect 165018 5366 165130 6646
rect 166200 5366 166312 6646
rect 167382 5366 167494 6646
rect 168564 5366 168676 6646
rect 169746 5366 169858 6646
rect 170928 5366 171040 6646
rect 172110 5366 172222 6646
rect 173292 5366 173404 6646
rect 174474 5366 174586 6646
rect 175656 5366 175768 6646
rect 176838 5366 176950 6646
rect 178020 5366 178132 6646
rect 179202 5366 179314 6646
rect 180384 5366 180496 6646
rect 181566 5366 181678 6646
rect 182748 5366 182860 6646
rect 183930 5366 184042 6646
rect 185112 5366 185224 6646
rect 186294 5366 186406 6646
rect 187476 5366 187588 6646
rect 188658 5366 188770 6646
rect 189840 5366 189952 6646
rect 191022 5366 191134 6646
rect 192204 5366 192316 6646
rect 193386 5366 193498 6646
rect 194568 5366 194680 6646
rect 195750 5366 195862 6646
rect 196932 5366 197044 6646
rect 198114 5366 198226 6646
rect 199296 5366 199408 6646
rect 200478 5366 200590 6646
rect 201660 5366 201772 6646
rect 202842 5366 202954 6646
rect 204024 5366 204136 6646
rect 205206 5366 205318 6646
rect 206388 5366 206500 6646
rect 207570 5366 207682 6646
rect 208752 5366 208864 6646
rect 209934 5366 210046 6646
rect 211116 5366 211228 6646
rect 212298 5366 212410 6646
rect 213480 5366 213592 6646
rect 214662 5366 214774 6646
rect 215844 5366 215956 6646
rect 217026 5366 217138 6646
rect 218208 5366 218320 6646
rect 219390 5366 219502 6646
rect 220572 5366 220684 6646
rect 221754 5366 221866 6646
rect 222936 5366 223048 6646
rect 224118 5366 224230 6646
rect 225300 5366 225412 6646
rect 226482 5366 226594 6646
rect 227664 5366 227776 6646
rect 228846 5366 228958 6646
rect 230028 5366 230140 6646
rect 231210 5366 231322 6646
rect 232392 5366 232504 6646
rect 233574 5366 233686 6646
rect 234756 5366 234868 6646
rect 235938 5366 236050 6646
rect 237120 5366 237232 6646
rect 238302 5366 238414 6646
rect 239484 5366 239596 6646
rect 240666 5366 240778 6646
rect 241848 5366 241960 6646
rect 243030 5366 243142 6646
rect 244212 5366 244324 6646
rect 245394 5366 245506 6646
rect 246576 5366 246688 6646
rect 247758 5366 247870 6646
rect 248940 5366 249052 6646
rect 250122 5366 250234 6646
rect 251304 5366 251416 6646
rect 252486 5366 252598 6646
rect 253668 5366 253780 6646
rect 254850 5366 254962 6646
rect 256032 5366 256144 6646
rect 257214 5366 257326 6646
rect 258396 5366 258508 6646
rect 259578 5366 259690 6646
rect 260760 5366 260872 6646
rect 261942 5366 262054 6646
rect 263124 5366 263236 6646
rect 264306 5366 264418 6646
rect 265488 5366 265600 6646
rect 266670 5366 266782 6646
rect 267852 5366 267964 6646
rect 269034 5366 269146 6646
rect 270216 5366 270328 6646
rect 271398 5366 271510 6646
rect 272580 5366 272692 6646
rect 273762 5366 273874 6646
rect 274944 5366 275056 6646
rect 276126 5366 276238 6646
rect 277308 5366 277420 6646
rect 278490 5366 278602 6646
rect 279672 5366 279784 6646
rect 280854 5366 280966 6646
rect 282036 5366 282148 6646
rect 283218 5366 283330 6646
rect 284400 5366 284512 6646
rect 285582 5366 285694 6646
rect 286764 5366 286876 6646
rect 287946 5366 288058 6646
rect 289128 5366 289240 6646
rect 290310 5366 290422 6646
rect 291492 5366 291604 6646
rect 292674 5366 292786 6646
rect 293856 5366 293968 6646
rect 295038 5366 295150 6646
rect 296220 5366 296332 6646
rect 297402 5366 297514 6646
rect 298584 5366 298696 6646
rect 299766 5366 299878 6646
rect 300948 5366 301060 6646
rect 302130 5366 302242 6646
rect 303312 5366 303424 6646
rect 304494 5366 304606 6646
rect 305676 5366 305788 6646
rect 306858 5366 306970 6646
rect 308040 5366 308152 6646
rect 309222 5366 309334 6646
rect 310404 5366 310516 6646
rect 311586 5366 311698 6646
rect 312768 5366 312880 6646
rect 313950 5366 314062 6646
rect 315132 5366 315244 6646
rect 316314 5366 316426 6646
rect 317496 5366 317608 6646
rect 318678 5366 318790 6646
rect 319860 5366 319972 6646
rect 321042 5366 321154 6646
rect 322224 5366 322336 6646
rect 323406 5366 323518 6646
rect 324588 5366 324700 6646
rect 325770 5366 325882 6646
rect 326952 5366 327064 6646
rect 328134 5366 328246 6646
rect 329316 5366 329428 6646
rect 330498 5366 330610 6646
rect 331680 5366 331792 6646
rect 332862 5366 332974 6646
rect 334044 5366 334156 6646
rect 335226 5366 335338 6646
rect 336408 5366 336520 6646
rect 337590 5366 337702 6646
rect 338772 5366 338884 6646
rect 339954 5366 340066 6646
rect 341136 5366 341248 6646
rect 342318 5366 342430 6646
rect 343500 5366 343612 6646
rect 344682 5366 344794 6646
rect 345864 5366 345976 6646
rect 347046 5366 347158 6646
rect 348228 5366 348340 6646
rect 349410 5366 349522 6646
rect 350592 5366 350704 6646
rect 351774 5366 351886 6646
rect 352956 5366 353068 6646
rect 354138 5366 354250 6646
rect 355320 5366 355432 6646
rect 356502 5366 356614 6646
rect 357684 5366 357796 6646
rect 358866 5366 358978 6646
rect 360048 5366 360160 6646
rect 361230 5366 361342 6646
rect 362412 5366 362524 6646
rect 363594 5366 363706 6646
rect 364776 5366 364888 6646
rect 365958 5366 366070 6646
rect 367140 5366 367252 6646
rect 368322 5366 368434 6646
rect 369504 5366 369616 6646
rect 370686 5366 370798 6646
rect 371868 5366 371980 6646
rect 373050 5366 373162 6646
rect 374232 5366 374344 6646
rect 375414 5366 375526 6646
rect 376596 5366 376708 6646
rect 377778 5366 377890 6646
rect 378960 5366 379072 6646
rect 380142 5366 380254 6646
rect 381324 5366 381436 6646
rect 382506 5366 382618 6646
rect 383688 5366 383800 6646
rect 384870 5366 384982 6646
rect 386052 5366 386164 6646
rect 387234 5366 387346 6646
rect 388416 5366 388528 6646
rect 389598 5366 389710 6646
rect 390780 5366 390892 6646
rect 391962 5366 392074 6646
rect 393144 5366 393256 6646
rect 394326 5366 394438 6646
rect 395508 5366 395620 6646
rect 396690 5366 396802 6646
rect 397872 5366 397984 6646
rect 399054 5366 399166 6646
rect 400236 5366 400348 6646
rect 401418 5366 401530 6646
rect 402600 5366 402712 6646
rect 403782 5366 403894 6646
rect 404964 5366 405076 6646
rect 406146 5366 406258 6646
rect 407328 5366 407440 6646
rect 408510 5366 408622 6646
rect 409692 5366 409804 6646
rect 410874 5366 410986 6646
rect 412056 5366 412168 6646
rect 413238 5366 413350 6646
rect 414420 5366 414532 6646
rect 415602 5366 415714 6646
rect 416784 5366 416896 6646
rect 417966 5366 418078 6646
rect 419148 5366 419260 6646
rect 420330 5366 420442 6646
rect 421512 5366 421624 6646
rect 422694 5366 422806 6646
rect 423876 5366 423988 6646
rect 425058 5366 425170 6646
rect 426240 5366 426352 6646
rect 427422 5366 427534 6646
rect 428604 5366 428716 6646
rect 429786 5366 429898 6646
rect 430968 5366 431080 6646
rect 432150 5366 432262 6646
rect 433332 5366 433444 6646
rect 434514 5366 434626 6646
rect 435696 5366 435808 6646
rect 436878 5366 436990 6646
rect 438060 5366 438172 6646
rect 439242 5366 439354 6646
rect 440424 5366 440536 6646
rect 441606 5366 441718 6646
rect 442788 5366 442900 6646
rect 443970 5366 444082 6646
rect 445152 5366 445264 6646
rect 446334 5366 446446 6646
rect 447516 5366 447628 6646
rect 448698 5366 448810 6646
rect 449880 5366 449992 6646
rect 451062 5366 451174 6646
rect 452244 5366 452356 6646
rect 453426 5366 453538 6646
rect 454608 5366 454720 6646
rect 455790 5366 455902 6646
rect 456972 5366 457084 6646
rect 458154 5366 458266 6646
rect 459336 5366 459448 6646
rect 460518 5366 460630 6646
rect 461700 5366 461812 6646
rect 462882 5366 462994 6646
rect 464064 5366 464176 6646
rect 465246 5366 465358 6646
rect 466428 5366 466540 6646
rect 467610 5366 467722 6646
rect 468792 5366 468904 6646
rect 469974 5366 470086 6646
rect 471156 5366 471268 6646
rect 472338 5366 472450 6646
rect 473520 5366 473632 6646
rect 474702 5366 474814 6646
rect 475884 5366 475996 6646
rect 477066 5366 477178 6646
rect 478248 5366 478360 6646
rect 479430 5366 479542 6646
rect 480612 5366 480724 6646
rect 481794 5366 481906 6646
rect 482976 5366 483088 6646
rect 484158 5366 484270 6646
rect 485340 5366 485452 6646
rect 486522 5366 486634 6646
rect 487704 5366 487816 6646
rect 488886 5366 488998 6646
rect 490068 5366 490180 6646
rect 491250 5366 491362 6646
rect 492432 5366 492544 6646
rect 493614 5366 493726 6646
rect 494796 5366 494908 6646
rect 495978 5366 496090 6646
rect 497160 5366 497272 6646
rect 498342 5366 498454 6646
rect 499524 5366 499636 6646
rect 500706 5366 500818 6646
rect 501888 5366 502000 6646
rect 503070 5366 503182 6646
rect 504252 5366 504364 6646
rect 505434 5366 505546 6646
rect 506616 5366 506728 6646
rect 507798 5366 507910 6646
rect 508980 5366 509092 6646
rect 510162 5366 510274 6646
rect 511344 5366 511456 6646
rect 512526 5366 512638 6646
rect 513708 5366 513820 6646
rect 514890 5366 515002 6646
rect 516072 5366 516184 6646
rect 517254 5366 517366 6646
rect 518436 5366 518548 6646
rect 519618 5366 519730 6646
rect 520800 5366 520912 6646
rect 521982 5366 522094 6646
rect 523164 5366 523276 6646
rect 524346 5366 524458 6646
rect 525528 5366 525640 6646
rect 526710 5366 526822 6646
rect 527892 5366 528004 6646
rect 529074 5366 529186 6646
rect 530256 5366 530368 6646
rect 531438 5366 531550 6646
rect 532620 5366 532732 6646
rect 533802 5366 533914 6646
rect 534984 5366 535096 6646
rect 536166 5366 536278 6646
rect 537348 5366 537460 6646
rect 538530 5366 538642 6646
rect 539712 5366 539824 6646
rect 540894 5366 541006 6646
rect 542076 5366 542188 6646
rect 543258 5366 543370 6646
rect 544440 5366 544552 6646
rect 545622 5366 545734 6646
rect 546804 5366 546916 6646
rect 547986 5366 548098 6646
rect 549168 5366 549280 6646
rect 550350 5366 550462 6646
rect 551532 5366 551644 6646
rect 552714 5366 552826 6646
rect 553896 5366 554008 6646
rect 555078 5366 555190 6646
rect 556260 5366 556372 6646
rect 557442 5366 557554 6646
rect 558624 5366 558736 6646
rect 559806 5366 559918 6646
rect 560988 5366 561100 6646
rect 562170 5366 562282 6646
rect 563352 5366 563464 6646
rect 564534 5366 564646 6646
rect 565716 5366 565828 6646
rect 566898 5366 567010 6646
rect 568080 5366 568192 6646
rect 569262 5366 569374 6646
rect 570444 5366 570556 6646
rect 571626 5366 571738 6646
rect 572808 5366 572920 6646
rect 573990 5366 574102 6646
rect 575172 5366 575284 6646
rect 576354 5366 576466 6646
<< via2 >>
rect 350642 634223 352492 635565
<< metal3 >>
rect 9298 708466 14298 710166
rect 61298 708466 66298 710166
rect 113298 708466 118298 710166
rect 158698 708466 163698 710166
rect 163998 696769 166198 710166
rect -6896 686408 -5196 691408
rect 163998 689930 166198 690493
rect 166498 696769 168698 710166
rect 168998 708466 173998 710166
rect 210398 708466 215398 710166
rect 166498 689930 168698 690493
rect 215698 696802 217898 710166
rect 215698 690079 217898 690526
rect 218198 696802 220398 710166
rect 220698 708466 225698 710166
rect 218198 690079 220398 690526
rect 312098 655663 317098 710166
rect 317398 696784 319598 710166
rect 319898 700458 322098 710166
rect 322398 700458 327398 710166
rect 406498 708466 411498 710166
rect 458498 708466 463498 710166
rect 319898 698258 327398 700458
rect 317398 690204 319598 690510
rect -6896 650008 -5236 654808
rect 312098 649149 317098 649906
rect 322398 655663 327398 698258
rect 322398 649149 327398 649906
rect 503698 696730 508498 710166
rect -6896 640008 -5236 644808
rect 503698 643764 508498 690498
rect 503698 637282 508498 637946
rect 513698 696730 518498 710166
rect 559698 708466 564698 710166
rect 513698 643764 518498 690498
rect 575404 684150 577104 689150
rect 553154 645950 553670 650750
rect 559846 645950 577104 650750
rect 513698 637282 518498 637946
rect 553154 635950 553670 640750
rect 559846 635950 577104 640750
rect 350574 635565 352546 635623
rect 350574 634223 350642 635565
rect 352492 634223 352546 635565
rect 350574 634156 352546 634223
rect 333064 626460 338764 626529
rect 364203 626468 526713 626537
rect -6896 565608 -5236 570408
rect -6896 555608 -5236 560408
rect 333064 517808 333176 626460
rect 334837 625740 334843 625850
rect 334953 625803 334959 625850
rect 526193 625811 526199 625813
rect 334953 625743 338764 625803
rect 364203 625751 526199 625811
rect 526193 625749 526199 625751
rect 526263 625749 526269 625813
rect 334953 625740 334959 625743
rect 526209 625446 526215 625448
rect -7696 517696 333176 517808
rect 334071 625378 338764 625438
rect 364203 625386 526215 625446
rect 526209 625384 526215 625386
rect 526279 625384 526285 625448
rect -7696 516514 -6416 516626
rect -7696 515332 -6416 515444
rect -7696 514150 -6416 514262
rect -7696 512968 -6416 513080
rect -7696 511786 -6416 511898
rect -7696 474474 -6416 474586
rect -7696 473292 -6416 473404
rect -7696 472110 -6416 472222
rect -7696 470928 -6416 471040
rect 334071 469858 334183 625378
rect -7696 469746 334183 469858
rect 334842 624798 334954 624804
rect -7696 468564 6998 468676
rect 10668 468564 10815 468676
rect -7696 431252 -6416 431364
rect -7696 430070 -6416 430182
rect -7696 428888 -6416 429000
rect -7696 427706 -6416 427818
rect 334842 426636 334954 624686
rect -7696 426524 334954 426636
rect -7696 425342 6991 425454
rect 10703 425342 10798 425454
rect 526601 411574 526713 626468
rect 526998 625813 527062 625819
rect 527062 625751 532710 625811
rect 526998 625743 527062 625749
rect 527008 625448 527072 625454
rect 527072 625386 530592 625446
rect 527008 625378 527072 625384
rect 530480 460724 530592 625386
rect 532598 505146 532710 625751
rect 576624 595638 577904 595750
rect 576624 594456 577904 594568
rect 576624 593274 577904 593386
rect 576624 592092 577904 592204
rect 576624 590910 577904 591022
rect 576624 589728 577904 589840
rect 548556 556728 549333 561528
rect 555450 556728 577104 561528
rect 548556 546728 549333 551528
rect 555450 546728 577104 551528
rect 566475 506216 566652 506328
rect 569847 506216 577904 506328
rect 532598 505034 577904 505146
rect 576624 503852 577904 503964
rect 576624 502670 577904 502782
rect 576624 501488 577904 501600
rect 576624 500306 577904 500418
rect 566509 461794 566660 461906
rect 569835 461794 577904 461906
rect 530480 460612 577904 460724
rect 576624 459430 577904 459542
rect 576624 458248 577904 458360
rect 576624 457066 577904 457178
rect 576624 455884 577904 455996
rect 576624 417372 577904 417484
rect 576624 416190 577904 416302
rect 576624 415008 577904 415120
rect 576624 413826 577904 413938
rect 576624 412644 577904 412756
rect 526601 411462 577904 411574
rect -7696 388030 -6416 388142
rect -7696 386848 -6416 386960
rect -7696 385666 -6416 385778
rect -7696 384484 -6416 384596
rect -7696 383302 -6416 383414
rect -7696 382120 -6416 382232
rect 576624 370950 577904 371062
rect 576624 369768 577904 369880
rect 576624 368586 577904 368698
rect 576624 367404 577904 367516
rect 576624 366222 577904 366334
rect 576624 365040 577904 365152
rect -7696 344808 -6416 344920
rect -7696 343626 -6416 343738
rect -7696 342444 -6416 342556
rect -7696 341262 -6416 341374
rect -7696 340080 -6416 340192
rect -7696 338898 -6416 339010
rect 576624 325728 577904 325840
rect 576624 324546 577904 324658
rect 576624 323364 577904 323476
rect 576624 322182 577904 322294
rect 576624 321000 577904 321112
rect 576624 319818 577904 319930
rect -7696 301586 -6416 301698
rect -7696 300404 -6416 300516
rect -7696 299222 -6416 299334
rect -7696 298040 -6416 298152
rect -7696 296858 -6416 296970
rect -7696 295676 -6416 295788
rect 576624 281306 577904 281418
rect 576624 280124 577904 280236
rect 576624 278942 577904 279054
rect 576624 277760 577904 277872
rect 576624 276578 577904 276690
rect 576624 275396 577904 275508
rect -7696 258564 -6416 258676
rect -7696 257382 -6416 257494
rect -7696 256200 -6416 256312
rect -7696 255018 -6416 255130
rect -7696 253836 -6416 253948
rect -7696 252654 -6416 252766
rect 575444 241396 577104 246196
rect 575444 231396 577104 236196
rect -6896 221054 -5236 225854
rect -6896 211054 -5236 215854
rect 6510 197596 7095 202396
rect 10531 197596 566709 202396
rect 569733 197596 577104 202396
rect 575444 187596 577104 192396
rect -6896 179054 -5236 183854
rect -6896 169054 -5236 173854
rect 575444 152996 577104 157796
rect 575444 142996 577104 147796
rect -7696 130942 -6416 131054
rect -7696 129760 -6416 129872
rect -7696 128578 -6416 128690
rect -7696 127396 -6416 127508
rect -7696 126214 -6416 126326
rect -7696 125032 -6416 125144
rect 576624 101284 577904 101396
rect 576624 100102 577904 100214
rect 576624 98920 577904 99032
rect 576624 97738 577904 97850
rect -7696 87720 -6416 87832
rect -7696 86538 -6416 86650
rect -7696 85356 -6416 85468
rect -7696 84174 -6416 84286
rect -7696 82992 -6416 83104
rect -7696 81810 -6416 81922
rect 576624 56626 577904 56738
rect 576624 55444 577904 55556
rect 576624 54262 577904 54374
rect 576624 53080 577904 53192
rect -7696 44498 -6416 44610
rect -7696 43316 -6416 43428
rect -7696 42134 -6416 42246
rect -7696 40952 -6416 41064
rect -7696 39770 -6416 39882
rect -7696 38588 -6416 38700
rect 576624 30168 577904 30280
rect 576624 28986 577904 29098
rect 576624 27804 577904 27916
rect 576624 26622 577904 26734
rect 576624 25440 577904 25552
rect 576624 24258 577904 24370
rect -7696 23076 -6416 23188
rect 576624 23076 577904 23188
rect -7696 21894 -6416 22006
rect 576624 21894 577904 22006
rect -7696 20712 -6416 20824
rect 576624 20712 577904 20824
rect -7696 19530 -6416 19642
rect 576624 19530 577904 19642
rect -7696 18348 -6416 18460
rect 576624 18348 577904 18460
rect -7696 17166 -6416 17278
rect 576624 17166 577904 17278
rect -7696 15984 -6416 16096
rect 576624 15984 577904 16096
rect -7696 14802 -6416 14914
rect 576624 14802 577904 14914
rect -7696 13620 -6416 13732
rect 576624 13620 577904 13732
rect -7696 12438 -6416 12550
rect 576624 12438 577904 12550
rect -7696 11256 -6416 11368
rect 576624 11256 577904 11368
rect -7696 10074 -6416 10186
rect 576624 10074 577904 10186
rect -7696 8892 -6416 9004
rect 576624 8892 577904 9004
rect -7696 7710 -6416 7822
rect 576624 7710 577904 7822
<< via3 >>
rect 163998 690493 166198 696769
rect 166498 690493 168698 696769
rect 215698 690526 217898 696802
rect 218198 690526 220398 696802
rect 317398 690510 319598 696784
rect 312098 649906 317098 655663
rect 322398 649906 327398 655663
rect 503698 690498 508498 696730
rect 503698 637946 508498 643764
rect 513698 690498 518498 696730
rect 553670 645950 559846 650750
rect 513698 637946 518498 643764
rect 553670 635950 559846 640750
rect 350642 634223 352492 635565
rect 334843 625740 334953 625850
rect 526199 625749 526263 625813
rect 526215 625384 526279 625448
rect 334842 624686 334954 624798
rect 6998 468564 10668 468676
rect 6991 425342 10703 425454
rect 526998 625749 527062 625813
rect 527008 625384 527072 625448
rect 549333 556728 555450 561528
rect 549333 546728 555450 551528
rect 566652 506216 569847 506328
rect 566660 461794 569835 461906
rect 7095 197596 10531 202396
rect 566709 197596 569733 202396
<< metal4 >>
rect 163732 696802 519266 696903
rect 163732 696769 215698 696802
rect 163732 690493 163998 696769
rect 166198 690493 166498 696769
rect 168698 690526 215698 696769
rect 217898 690526 218198 696802
rect 220398 696784 519266 696802
rect 220398 690526 317398 696784
rect 168698 690510 317398 690526
rect 319598 696730 519266 696784
rect 319598 690510 503698 696730
rect 168698 690498 503698 690510
rect 508498 690498 513698 696730
rect 518498 690498 519266 696730
rect 168698 690493 519266 690498
rect 163732 690349 519266 690493
rect 311434 656003 353077 656064
rect 311434 655663 350663 656003
rect 311434 649906 312098 655663
rect 317098 649906 322398 655663
rect 327398 649906 350663 655663
rect 311434 649560 350663 649906
rect 352418 649560 353077 656003
rect 311434 649510 353077 649560
rect 553529 650750 560083 651146
rect 553529 645950 553670 650750
rect 559846 645950 560083 650750
rect 349248 643764 518800 644064
rect 349248 637946 503698 643764
rect 508498 637946 513698 643764
rect 518498 637946 518800 643764
rect 349248 637510 518800 637946
rect 553529 640750 560083 645950
rect 350546 635565 352574 637510
rect 350546 634223 350642 635565
rect 352492 634223 352574 635565
rect 350546 626039 352574 634223
rect 553529 635950 553670 640750
rect 559846 635950 560083 640750
rect 334842 625850 334954 625851
rect 334842 625740 334843 625850
rect 334953 625740 334954 625850
rect 334842 624799 334954 625740
rect 349971 625639 352989 626039
rect 526198 625813 526264 625814
rect 526198 625749 526199 625813
rect 526263 625811 526264 625813
rect 526997 625813 527063 625814
rect 526997 625811 526998 625813
rect 526263 625751 526998 625811
rect 526263 625749 526264 625751
rect 526198 625748 526264 625749
rect 526997 625749 526998 625751
rect 527062 625749 527063 625813
rect 526997 625748 527063 625749
rect 526214 625448 526280 625449
rect 526214 625384 526215 625448
rect 526279 625446 526280 625448
rect 527007 625448 527073 625449
rect 527007 625446 527008 625448
rect 526279 625386 527008 625446
rect 526279 625384 526280 625386
rect 526214 625383 526280 625384
rect 527007 625384 527008 625386
rect 527072 625384 527073 625448
rect 527007 625383 527073 625384
rect 334841 624798 334955 624799
rect 334841 624686 334842 624798
rect 334954 624686 334955 624798
rect 334841 624685 334955 624686
rect 338877 619922 339932 625015
rect 345032 623995 346861 625022
rect 345032 621415 345132 623995
rect 346707 621415 346861 623995
rect 345032 621297 346861 621415
rect 356432 624001 358261 625050
rect 356432 621421 356516 624001
rect 358091 621421 358261 624001
rect 356432 621297 358261 621421
rect 362927 619922 364084 625025
rect 553529 619922 560083 635950
rect 338360 613368 560083 619922
rect 355762 607738 555717 607922
rect 355762 603397 356518 607738
rect 358096 603397 555717 607738
rect 355762 601368 555717 603397
rect 549163 561528 555717 601368
rect 549163 556728 549333 561528
rect 555450 556728 555717 561528
rect 549163 551528 555717 556728
rect 549163 546728 549333 551528
rect 555450 546728 555717 551528
rect 549163 546321 555717 546728
rect 566568 506328 569920 506639
rect 566568 506216 566652 506328
rect 569847 506216 569920 506328
rect 6918 468676 10788 468937
rect 6918 468564 6998 468676
rect 10668 468564 10788 468676
rect 6918 425454 10788 468564
rect 6918 425342 6991 425454
rect 10703 425342 10788 425454
rect 6918 233423 10788 425342
rect 566568 461906 569920 506216
rect 566568 461794 566660 461906
rect 569835 461794 569920 461906
rect 6915 202396 10792 233423
rect 6915 197596 7095 202396
rect 10531 197596 10792 202396
rect 6915 197264 10792 197596
rect 566568 202396 569920 461794
rect 566568 197596 566709 202396
rect 569733 197596 569920 202396
rect 566568 197357 569920 197596
<< via4 >>
rect 350663 649560 352418 656003
rect 345132 621415 346707 623995
rect 356516 621421 358091 624001
rect 356518 603397 358096 607738
<< metal5 >>
rect 350625 656003 352454 656157
rect 350625 649560 350663 656003
rect 352418 649560 352454 656003
rect 345022 623995 346851 624095
rect 345022 621415 345132 623995
rect 346707 621415 346851 623995
rect 345022 621066 346851 621415
rect 350625 621066 352454 649560
rect 345022 619237 352454 621066
rect 356422 624001 358251 624095
rect 356422 621421 356516 624001
rect 358091 621421 358251 624001
rect 356422 607738 358251 621421
rect 356422 603397 356518 607738
rect 358096 603397 358251 607738
rect 356422 603218 358251 603397
<< comment >>
rect -6996 710166 577204 710266
rect -6996 6166 -6896 710166
rect 577104 6166 577204 710166
rect -6996 6066 577204 6166
use user_analog_proj_example  user_analog_proj_example_0
timestamp 1620310959
transform 1 0 338772 0 -1 633280
box -59 -22 25476 8324
<< labels >>
flabel metal3 s 576624 275396 577904 275508 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -7696 388030 -6416 388142 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -7696 344808 -6416 344920 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -7696 301586 -6416 301698 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -7696 258564 -6416 258676 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -7696 130942 -6416 131054 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -7696 87720 -6416 87832 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -7696 44498 -6416 44610 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -7696 23076 -6416 23188 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 576624 319818 577904 319930 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 576624 365040 577904 365152 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 576624 411462 577904 411574 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 576624 455884 577904 455996 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 576624 500306 577904 500418 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 576624 589728 577904 589840 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -7696 517696 -6416 517808 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -7696 474474 -6416 474586 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -7696 431252 -6416 431364 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 576624 276578 577904 276690 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -7696 386848 -6416 386960 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -7696 343626 -6416 343738 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -7696 300404 -6416 300516 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -7696 257382 -6416 257494 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -7696 129760 -6416 129872 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -7696 86538 -6416 86650 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -7696 43316 -6416 43428 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -7696 21894 -6416 22006 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 576624 321000 577904 321112 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 576624 366222 577904 366334 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 576624 412644 577904 412756 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 576624 457066 577904 457178 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 576624 501488 577904 501600 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 576624 590910 577904 591022 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -7696 516514 -6416 516626 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -7696 473292 -6416 473404 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -7696 430070 -6416 430182 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 575404 684150 577104 689150 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s -6896 686408 -5196 691408 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 559698 708466 564698 710166 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 458498 708466 463498 710166 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 406498 708466 411498 710166 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 322398 708466 327398 710166 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 220698 708466 225698 710166 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 168998 708466 173998 710166 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 113298 708466 118298 710166 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 61298 708466 66298 710166 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 9298 708466 14298 710166 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 312098 708466 317098 710166 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 210398 708466 215398 710166 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 158698 708466 163698 710166 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 319898 708466 322098 710166 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 218198 708466 220398 710166 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 166498 708466 168698 710166 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 317398 708466 319598 710166 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 215698 708466 217898 710166 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 163998 708466 166198 710166 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 576624 8892 577904 9004 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 576624 415008 577904 415120 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 576624 459430 577904 459542 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 576624 503852 577904 503964 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 576624 593274 577904 593386 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -7696 514150 -6416 514262 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -7696 470928 -6416 471040 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -7696 427706 -6416 427818 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -7696 384484 -6416 384596 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -7696 341262 -6416 341374 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -7696 298040 -6416 298152 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 576624 13620 577904 13732 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -7696 255018 -6416 255130 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -7696 127396 -6416 127508 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -7696 84174 -6416 84286 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -7696 40952 -6416 41064 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -7696 19530 -6416 19642 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -7696 14802 -6416 14914 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -7696 10074 -6416 10186 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 576624 18348 577904 18460 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 576624 23076 577904 23188 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 576624 27804 577904 27916 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 576624 54262 577904 54374 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 576624 98920 577904 99032 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 576624 278942 577904 279054 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 576624 323364 577904 323476 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 576624 368586 577904 368698 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 576624 7710 577904 7822 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 576624 413826 577904 413938 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 576624 458248 577904 458360 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 576624 502670 577904 502782 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 576624 592092 577904 592204 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -7696 515332 -6416 515444 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -7696 472110 -6416 472222 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -7696 428888 -6416 429000 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -7696 385666 -6416 385778 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -7696 342444 -6416 342556 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -7696 299222 -6416 299334 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 576624 12438 577904 12550 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -7696 256200 -6416 256312 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -7696 128578 -6416 128690 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -7696 85356 -6416 85468 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -7696 42134 -6416 42246 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -7696 20712 -6416 20824 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -7696 15984 -6416 16096 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -7696 11256 -6416 11368 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 576624 17166 577904 17278 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 576624 21894 577904 22006 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 576624 26622 577904 26734 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 576624 53080 577904 53192 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 576624 97738 577904 97850 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 576624 277760 577904 277872 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 576624 322182 577904 322294 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 576624 367404 577904 367516 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 576624 11256 577904 11368 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 576624 417372 577904 417484 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 576624 461794 577904 461906 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 576624 506216 577904 506328 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 576624 595638 577904 595750 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -7696 511786 -6416 511898 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -7696 468564 -6416 468676 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -7696 425342 -6416 425454 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -7696 382120 -6416 382232 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -7696 338898 -6416 339010 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -7696 295676 -6416 295788 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 576624 15984 577904 16096 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -7696 252654 -6416 252766 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -7696 125032 -6416 125144 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -7696 81810 -6416 81922 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -7696 38588 -6416 38700 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -7696 17166 -6416 17278 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -7696 12438 -6416 12550 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -7696 7710 -6416 7822 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 576624 20712 577904 20824 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 576624 25440 577904 25552 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 576624 30168 577904 30280 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 576624 56626 577904 56738 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 576624 101284 577904 101396 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 576624 281306 577904 281418 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 576624 325728 577904 325840 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 576624 370950 577904 371062 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 576624 10074 577904 10186 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 576624 416190 577904 416302 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 576624 460612 577904 460724 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 576624 505034 577904 505146 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 576624 594456 577904 594568 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -7696 512968 -6416 513080 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -7696 469746 -6416 469858 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -7696 426524 -6416 426636 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -7696 383302 -6416 383414 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -7696 340080 -6416 340192 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -7696 296858 -6416 296970 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 576624 14802 577904 14914 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -7696 253836 -6416 253948 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -7696 126214 -6416 126326 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -7696 82992 -6416 83104 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -7696 39770 -6416 39882 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -7696 18348 -6416 18460 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -7696 13620 -6416 13732 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -7696 8892 -6416 9004 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 576624 19530 577904 19642 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 576624 24258 577904 24370 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 576624 28986 577904 29098 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 576624 55444 577904 55556 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 576624 100102 577904 100214 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 576624 280124 577904 280236 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 576624 324546 577904 324658 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 576624 369768 577904 369880 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 118920 5366 119032 6646 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 473520 5366 473632 6646 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 477066 5366 477178 6646 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 480612 5366 480724 6646 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 484158 5366 484270 6646 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 487704 5366 487816 6646 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 491250 5366 491362 6646 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 494796 5366 494908 6646 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 498342 5366 498454 6646 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 501888 5366 502000 6646 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 505434 5366 505546 6646 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 154380 5366 154492 6646 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 508980 5366 509092 6646 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 512526 5366 512638 6646 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 516072 5366 516184 6646 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 519618 5366 519730 6646 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 523164 5366 523276 6646 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 526710 5366 526822 6646 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 530256 5366 530368 6646 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 533802 5366 533914 6646 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 537348 5366 537460 6646 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 540894 5366 541006 6646 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 157926 5366 158038 6646 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 544440 5366 544552 6646 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 547986 5366 548098 6646 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 551532 5366 551644 6646 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 555078 5366 555190 6646 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 558624 5366 558736 6646 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 562170 5366 562282 6646 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 565716 5366 565828 6646 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 569262 5366 569374 6646 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 161472 5366 161584 6646 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 165018 5366 165130 6646 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 168564 5366 168676 6646 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 172110 5366 172222 6646 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 175656 5366 175768 6646 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 179202 5366 179314 6646 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 182748 5366 182860 6646 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 186294 5366 186406 6646 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 122466 5366 122578 6646 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 189840 5366 189952 6646 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 193386 5366 193498 6646 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 196932 5366 197044 6646 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 200478 5366 200590 6646 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 204024 5366 204136 6646 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 207570 5366 207682 6646 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 211116 5366 211228 6646 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 214662 5366 214774 6646 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 218208 5366 218320 6646 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 221754 5366 221866 6646 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 126012 5366 126124 6646 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 225300 5366 225412 6646 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 228846 5366 228958 6646 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 232392 5366 232504 6646 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 235938 5366 236050 6646 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 239484 5366 239596 6646 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 243030 5366 243142 6646 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 246576 5366 246688 6646 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 250122 5366 250234 6646 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 253668 5366 253780 6646 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 257214 5366 257326 6646 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 129558 5366 129670 6646 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 260760 5366 260872 6646 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 264306 5366 264418 6646 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 267852 5366 267964 6646 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 271398 5366 271510 6646 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 274944 5366 275056 6646 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 278490 5366 278602 6646 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 282036 5366 282148 6646 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 285582 5366 285694 6646 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 289128 5366 289240 6646 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 292674 5366 292786 6646 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 133104 5366 133216 6646 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 296220 5366 296332 6646 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 299766 5366 299878 6646 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 303312 5366 303424 6646 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 306858 5366 306970 6646 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 310404 5366 310516 6646 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 313950 5366 314062 6646 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 317496 5366 317608 6646 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 321042 5366 321154 6646 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 324588 5366 324700 6646 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 328134 5366 328246 6646 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 136650 5366 136762 6646 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 331680 5366 331792 6646 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 335226 5366 335338 6646 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 338772 5366 338884 6646 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 342318 5366 342430 6646 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 345864 5366 345976 6646 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 349410 5366 349522 6646 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 352956 5366 353068 6646 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 356502 5366 356614 6646 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 360048 5366 360160 6646 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 363594 5366 363706 6646 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 140196 5366 140308 6646 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 367140 5366 367252 6646 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 370686 5366 370798 6646 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 374232 5366 374344 6646 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 377778 5366 377890 6646 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 381324 5366 381436 6646 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 384870 5366 384982 6646 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 388416 5366 388528 6646 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 391962 5366 392074 6646 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 395508 5366 395620 6646 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 399054 5366 399166 6646 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 143742 5366 143854 6646 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 402600 5366 402712 6646 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 406146 5366 406258 6646 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 409692 5366 409804 6646 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 413238 5366 413350 6646 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 416784 5366 416896 6646 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 420330 5366 420442 6646 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 423876 5366 423988 6646 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 427422 5366 427534 6646 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 430968 5366 431080 6646 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 434514 5366 434626 6646 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 147288 5366 147400 6646 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 438060 5366 438172 6646 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 441606 5366 441718 6646 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 445152 5366 445264 6646 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 448698 5366 448810 6646 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 452244 5366 452356 6646 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 455790 5366 455902 6646 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 459336 5366 459448 6646 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 462882 5366 462994 6646 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 466428 5366 466540 6646 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 469974 5366 470086 6646 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 150834 5366 150946 6646 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 120102 5366 120214 6646 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 474702 5366 474814 6646 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 478248 5366 478360 6646 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 481794 5366 481906 6646 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 485340 5366 485452 6646 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 488886 5366 488998 6646 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 492432 5366 492544 6646 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 495978 5366 496090 6646 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 499524 5366 499636 6646 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 503070 5366 503182 6646 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 506616 5366 506728 6646 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 155562 5366 155674 6646 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 510162 5366 510274 6646 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 513708 5366 513820 6646 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 517254 5366 517366 6646 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 520800 5366 520912 6646 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 524346 5366 524458 6646 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 527892 5366 528004 6646 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 531438 5366 531550 6646 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 534984 5366 535096 6646 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 538530 5366 538642 6646 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 542076 5366 542188 6646 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 159108 5366 159220 6646 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 545622 5366 545734 6646 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 549168 5366 549280 6646 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 552714 5366 552826 6646 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 556260 5366 556372 6646 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 559806 5366 559918 6646 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 563352 5366 563464 6646 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 566898 5366 567010 6646 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 570444 5366 570556 6646 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 162654 5366 162766 6646 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 166200 5366 166312 6646 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 169746 5366 169858 6646 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 173292 5366 173404 6646 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 176838 5366 176950 6646 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 180384 5366 180496 6646 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 183930 5366 184042 6646 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 187476 5366 187588 6646 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 123648 5366 123760 6646 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 191022 5366 191134 6646 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 194568 5366 194680 6646 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 198114 5366 198226 6646 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 201660 5366 201772 6646 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 205206 5366 205318 6646 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 208752 5366 208864 6646 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 212298 5366 212410 6646 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 215844 5366 215956 6646 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 219390 5366 219502 6646 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 222936 5366 223048 6646 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 127194 5366 127306 6646 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 226482 5366 226594 6646 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 230028 5366 230140 6646 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 233574 5366 233686 6646 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 237120 5366 237232 6646 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 240666 5366 240778 6646 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 244212 5366 244324 6646 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 247758 5366 247870 6646 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 251304 5366 251416 6646 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 254850 5366 254962 6646 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 258396 5366 258508 6646 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 130740 5366 130852 6646 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 261942 5366 262054 6646 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 265488 5366 265600 6646 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 269034 5366 269146 6646 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 272580 5366 272692 6646 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 276126 5366 276238 6646 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 279672 5366 279784 6646 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 283218 5366 283330 6646 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 286764 5366 286876 6646 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 290310 5366 290422 6646 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 293856 5366 293968 6646 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 134286 5366 134398 6646 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 297402 5366 297514 6646 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 300948 5366 301060 6646 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 304494 5366 304606 6646 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 308040 5366 308152 6646 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 311586 5366 311698 6646 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 315132 5366 315244 6646 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 318678 5366 318790 6646 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 322224 5366 322336 6646 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 325770 5366 325882 6646 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 329316 5366 329428 6646 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 137832 5366 137944 6646 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 332862 5366 332974 6646 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 336408 5366 336520 6646 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 339954 5366 340066 6646 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 343500 5366 343612 6646 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 347046 5366 347158 6646 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 350592 5366 350704 6646 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 354138 5366 354250 6646 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 357684 5366 357796 6646 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 361230 5366 361342 6646 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 364776 5366 364888 6646 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 141378 5366 141490 6646 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 368322 5366 368434 6646 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 371868 5366 371980 6646 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 375414 5366 375526 6646 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 378960 5366 379072 6646 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 382506 5366 382618 6646 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 386052 5366 386164 6646 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 389598 5366 389710 6646 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 393144 5366 393256 6646 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 396690 5366 396802 6646 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 400236 5366 400348 6646 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 144924 5366 145036 6646 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 403782 5366 403894 6646 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 407328 5366 407440 6646 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 410874 5366 410986 6646 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 414420 5366 414532 6646 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 417966 5366 418078 6646 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 421512 5366 421624 6646 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 425058 5366 425170 6646 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 428604 5366 428716 6646 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 432150 5366 432262 6646 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 435696 5366 435808 6646 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 148470 5366 148582 6646 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 439242 5366 439354 6646 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 442788 5366 442900 6646 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 446334 5366 446446 6646 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 449880 5366 449992 6646 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 453426 5366 453538 6646 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 456972 5366 457084 6646 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 460518 5366 460630 6646 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 464064 5366 464176 6646 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 467610 5366 467722 6646 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 471156 5366 471268 6646 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 152016 5366 152128 6646 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 121284 5366 121396 6646 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 475884 5366 475996 6646 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 479430 5366 479542 6646 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 482976 5366 483088 6646 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 486522 5366 486634 6646 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 490068 5366 490180 6646 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 493614 5366 493726 6646 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 497160 5366 497272 6646 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 500706 5366 500818 6646 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 504252 5366 504364 6646 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 507798 5366 507910 6646 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 156744 5366 156856 6646 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 511344 5366 511456 6646 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 514890 5366 515002 6646 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 518436 5366 518548 6646 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 521982 5366 522094 6646 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 525528 5366 525640 6646 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 529074 5366 529186 6646 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 532620 5366 532732 6646 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 536166 5366 536278 6646 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 539712 5366 539824 6646 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 543258 5366 543370 6646 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 160290 5366 160402 6646 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 546804 5366 546916 6646 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 550350 5366 550462 6646 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 553896 5366 554008 6646 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 557442 5366 557554 6646 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 560988 5366 561100 6646 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 564534 5366 564646 6646 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 568080 5366 568192 6646 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 571626 5366 571738 6646 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 163836 5366 163948 6646 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 167382 5366 167494 6646 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 170928 5366 171040 6646 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 174474 5366 174586 6646 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 178020 5366 178132 6646 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 181566 5366 181678 6646 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 185112 5366 185224 6646 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 188658 5366 188770 6646 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 124830 5366 124942 6646 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 192204 5366 192316 6646 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 195750 5366 195862 6646 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 199296 5366 199408 6646 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 202842 5366 202954 6646 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 206388 5366 206500 6646 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 209934 5366 210046 6646 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 213480 5366 213592 6646 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 217026 5366 217138 6646 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 220572 5366 220684 6646 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 224118 5366 224230 6646 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 128376 5366 128488 6646 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 227664 5366 227776 6646 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 231210 5366 231322 6646 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 234756 5366 234868 6646 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 238302 5366 238414 6646 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 241848 5366 241960 6646 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 245394 5366 245506 6646 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 248940 5366 249052 6646 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 252486 5366 252598 6646 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 256032 5366 256144 6646 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 259578 5366 259690 6646 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 131922 5366 132034 6646 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 263124 5366 263236 6646 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 266670 5366 266782 6646 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 270216 5366 270328 6646 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 273762 5366 273874 6646 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 277308 5366 277420 6646 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 280854 5366 280966 6646 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 284400 5366 284512 6646 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 287946 5366 288058 6646 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 291492 5366 291604 6646 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 295038 5366 295150 6646 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 135468 5366 135580 6646 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 298584 5366 298696 6646 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 302130 5366 302242 6646 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 305676 5366 305788 6646 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 309222 5366 309334 6646 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 312768 5366 312880 6646 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 316314 5366 316426 6646 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 319860 5366 319972 6646 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 323406 5366 323518 6646 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 326952 5366 327064 6646 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 330498 5366 330610 6646 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 139014 5366 139126 6646 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 334044 5366 334156 6646 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 337590 5366 337702 6646 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 341136 5366 341248 6646 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 344682 5366 344794 6646 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 348228 5366 348340 6646 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 351774 5366 351886 6646 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 355320 5366 355432 6646 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 358866 5366 358978 6646 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 362412 5366 362524 6646 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 365958 5366 366070 6646 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 142560 5366 142672 6646 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 369504 5366 369616 6646 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 373050 5366 373162 6646 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 376596 5366 376708 6646 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 380142 5366 380254 6646 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 383688 5366 383800 6646 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 387234 5366 387346 6646 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 390780 5366 390892 6646 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 394326 5366 394438 6646 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 397872 5366 397984 6646 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 401418 5366 401530 6646 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 146106 5366 146218 6646 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 404964 5366 405076 6646 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 408510 5366 408622 6646 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 412056 5366 412168 6646 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 415602 5366 415714 6646 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 419148 5366 419260 6646 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 422694 5366 422806 6646 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 426240 5366 426352 6646 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 429786 5366 429898 6646 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 433332 5366 433444 6646 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 436878 5366 436990 6646 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 149652 5366 149764 6646 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 440424 5366 440536 6646 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 443970 5366 444082 6646 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 447516 5366 447628 6646 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 451062 5366 451174 6646 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 454608 5366 454720 6646 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 458154 5366 458266 6646 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 461700 5366 461812 6646 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 465246 5366 465358 6646 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 468792 5366 468904 6646 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 472338 5366 472450 6646 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 153198 5366 153310 6646 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 572808 5366 572920 6646 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 573990 5366 574102 6646 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 575172 5366 575284 6646 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 576354 5366 576466 6646 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 575444 645950 577104 650750 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 575444 635950 577104 640750 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s -6896 650008 -5236 654808 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s -6896 640008 -5236 644808 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 575444 546728 577104 551528 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 575444 556728 577104 561528 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 575444 241396 577104 246196 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 575444 231396 577104 236196 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s -6896 211054 -5236 215854 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s -6896 221054 -5236 225854 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 513698 708506 518498 710166 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 503698 708506 508498 710166 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 575444 152996 577104 157796 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 575444 142996 577104 147796 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s -6896 565608 -5236 570408 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s -6896 555608 -5236 560408 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 575444 197596 577104 202396 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 575444 187596 577104 192396 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s -6896 179054 -5236 183854 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s -6896 169054 -5236 173854 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s -6372 5366 -6260 6646 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s -5190 5366 -5078 6646 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s -4008 5366 -3896 6646 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 720 5366 832 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 40908 5366 41020 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 44454 5366 44566 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 48000 5366 48112 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 51546 5366 51658 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 55092 5366 55204 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 58638 5366 58750 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 62184 5366 62296 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 65730 5366 65842 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 69276 5366 69388 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 72822 5366 72934 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 5448 5366 5560 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 76368 5366 76480 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 79914 5366 80026 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 83460 5366 83572 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 87006 5366 87118 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 90552 5366 90664 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 94098 5366 94210 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 97644 5366 97756 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 101190 5366 101302 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 104736 5366 104848 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 108282 5366 108394 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 10176 5366 10288 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 111828 5366 111940 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 115374 5366 115486 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 14904 5366 15016 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 19632 5366 19744 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 23178 5366 23290 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 26724 5366 26836 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 30270 5366 30382 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 33816 5366 33928 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 37362 5366 37474 6646 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s -2826 5366 -2714 6646 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 1902 5366 2014 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 42090 5366 42202 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 45636 5366 45748 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 49182 5366 49294 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 52728 5366 52840 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 56274 5366 56386 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 59820 5366 59932 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 63366 5366 63478 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 66912 5366 67024 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 70458 5366 70570 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 74004 5366 74116 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 6630 5366 6742 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 77550 5366 77662 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 81096 5366 81208 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 84642 5366 84754 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 88188 5366 88300 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 91734 5366 91846 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 95280 5366 95392 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 98826 5366 98938 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 102372 5366 102484 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 105918 5366 106030 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 109464 5366 109576 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 11358 5366 11470 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 113010 5366 113122 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 116556 5366 116668 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 16086 5366 16198 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 20814 5366 20926 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 24360 5366 24472 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 27906 5366 28018 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 31452 5366 31564 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 34998 5366 35110 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 38544 5366 38656 6646 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 3084 5366 3196 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 43272 5366 43384 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 46818 5366 46930 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 50364 5366 50476 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 53910 5366 54022 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 57456 5366 57568 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 61002 5366 61114 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 64548 5366 64660 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 68094 5366 68206 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 71640 5366 71752 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 75186 5366 75298 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 7812 5366 7924 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 78732 5366 78844 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 82278 5366 82390 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 85824 5366 85936 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 89370 5366 89482 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 92916 5366 93028 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 96462 5366 96574 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 100008 5366 100120 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 103554 5366 103666 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 107100 5366 107212 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 110646 5366 110758 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 12540 5366 12652 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 114192 5366 114304 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 117738 5366 117850 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 17268 5366 17380 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 21996 5366 22108 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 25542 5366 25654 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 29088 5366 29200 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 32634 5366 32746 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 36180 5366 36292 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 39726 5366 39838 6646 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 4266 5366 4378 6646 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 8994 5366 9106 6646 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 13722 5366 13834 6646 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 18450 5366 18562 6646 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s -1644 5366 -1532 6646 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s -462 5366 -350 6646 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 565256 646308 573324 650316 0 FreeSans 16000 0 0 0 VCCD1
flabel metal3 560142 557126 570406 560712 0 FreeSans 16000 0 0 0 VDDA1
flabel metal3 504294 671062 508066 682438 0 FreeSans 16000 90 0 0 VSSA1
flabel metal3 554807 198095 564825 202025 0 FreeSans 16000 0 0 0 VSSD1
<< end >>
