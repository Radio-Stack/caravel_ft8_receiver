magic
tech sky130A
magscale 1 2
timestamp 1619730755
<< error_s >>
rect 347036 623411 347056 623429
rect 361194 623403 361214 623421
rect 346970 623345 346990 623363
rect 361128 623337 361148 623355
<< metal2 >>
rect 19384 703508 19496 704948
rect 58300 703508 58412 704948
rect 97216 703508 97328 704948
rect 136132 703508 136244 704948
rect 175048 703508 175160 704948
rect 214056 703508 214168 704948
rect 252972 703508 253084 704948
rect 291888 703578 292000 704948
rect 330804 703508 330916 704948
rect 369720 704106 369832 704948
rect 365888 703508 366000 703578
rect 351354 628628 351968 628750
rect 351354 626932 351424 628628
rect 351850 626932 351968 628628
rect 351354 626848 351968 626932
rect 351503 623888 351733 626848
rect 349528 623658 351733 623888
rect 369514 623880 369970 704106
rect 408728 703508 408840 704948
rect 447644 703508 447756 704948
rect 486560 703508 486672 704948
rect 525476 703508 525588 704948
rect 564392 703508 564504 704948
rect 371198 644874 373412 644898
rect 371198 644684 371240 644874
rect 372084 644868 373412 644874
rect 372084 644690 372762 644868
rect 373386 644690 373412 644868
rect 372084 644684 373412 644690
rect 371198 644650 373412 644684
rect 370616 641666 373926 641696
rect 370616 641480 370660 641666
rect 371192 641664 373926 641666
rect 371192 641496 373272 641664
rect 373888 641496 373926 641664
rect 371192 641480 373926 641496
rect 370616 641454 373926 641480
rect 370984 637098 373694 637128
rect 370984 636912 371028 637098
rect 371560 637096 373694 637098
rect 371560 636928 373040 637096
rect 373656 636928 373694 637096
rect 371560 636912 373694 636928
rect 370984 636886 373694 636912
rect 371518 625304 371728 625327
rect 371518 624430 371548 625304
rect 371696 624430 371728 625304
rect 372758 624652 372974 624670
rect 371518 624398 371728 624430
rect 371976 624650 372148 624652
rect 371976 624632 372192 624650
rect 363664 623650 369970 623880
rect 371544 622902 371716 624398
rect 371976 624060 372000 624632
rect 372174 624324 372192 624632
rect 372758 624324 372782 624652
rect 372174 624080 372782 624324
rect 372956 624080 372974 624652
rect 372174 624076 372974 624080
rect 372174 624060 372192 624076
rect 372758 624060 372974 624076
rect 371976 624040 372192 624060
rect 372764 624054 372974 624060
rect 371982 624034 372192 624040
rect 371544 622884 371760 622902
rect 371544 622312 371568 622884
rect 371742 622312 371760 622884
rect 371544 622292 371760 622312
rect 371550 622286 371760 622292
rect 524 -972 636 468
rect 1628 -972 1740 468
rect 2824 -972 2936 468
rect 4020 -972 4132 468
rect 5216 -972 5328 468
rect 6412 -972 6524 468
rect 7608 -972 7720 468
rect 8712 -972 8824 468
rect 9908 -972 10020 468
rect 11104 -972 11216 468
rect 12300 -972 12412 468
rect 13496 -972 13608 468
rect 14692 -972 14804 468
rect 15888 -972 16000 468
rect 16992 -972 17104 468
rect 18188 -972 18300 468
rect 19384 -972 19496 468
rect 20580 -972 20692 468
rect 21776 -972 21888 468
rect 22972 -972 23084 468
rect 24168 -972 24280 468
rect 25272 -972 25384 468
rect 26468 -972 26580 468
rect 27664 -972 27776 468
rect 28860 -972 28972 468
rect 30056 -972 30168 468
rect 31252 -972 31364 468
rect 32356 -972 32468 468
rect 33552 -972 33664 468
rect 34748 -972 34860 468
rect 35944 -972 36056 468
rect 37140 -972 37252 468
rect 38336 -972 38448 468
rect 39532 -972 39644 468
rect 40636 -972 40748 468
rect 41832 -972 41944 468
rect 43028 -972 43140 468
rect 44224 -972 44336 468
rect 45420 -972 45532 468
rect 46616 -972 46728 468
rect 47812 -972 47924 468
rect 48916 -972 49028 468
rect 50112 -972 50224 468
rect 51308 -972 51420 468
rect 52504 -972 52616 468
rect 53700 -972 53812 468
rect 54896 -972 55008 468
rect 56000 -972 56112 468
rect 57196 -972 57308 468
rect 58392 -972 58504 468
rect 59588 -972 59700 468
rect 60784 -972 60896 468
rect 61980 -972 62092 468
rect 63176 -972 63288 468
rect 64280 -972 64392 468
rect 65476 -972 65588 468
rect 66672 -972 66784 468
rect 67868 -972 67980 468
rect 69064 -972 69176 468
rect 70260 -972 70372 468
rect 71456 -972 71568 468
rect 72560 -972 72672 468
rect 73756 -972 73868 468
rect 74952 -972 75064 468
rect 76148 -972 76260 468
rect 77344 -972 77456 468
rect 78540 -972 78652 468
rect 79644 -972 79756 468
rect 80840 -972 80952 468
rect 82036 -972 82148 468
rect 83232 -972 83344 468
rect 84428 -972 84540 468
rect 85624 -972 85736 468
rect 86820 -972 86932 468
rect 87924 -972 88036 468
rect 89120 -972 89232 468
rect 90316 -972 90428 468
rect 91512 -972 91624 468
rect 92708 -972 92820 468
rect 93904 -972 94016 468
rect 95100 -972 95212 468
rect 96204 -972 96316 468
rect 97400 -972 97512 468
rect 98596 -972 98708 468
rect 99792 -972 99904 468
rect 100988 -972 101100 468
rect 102184 -972 102296 468
rect 103288 -972 103400 468
rect 104484 -972 104596 468
rect 105680 -972 105792 468
rect 106876 -972 106988 468
rect 108072 -972 108184 468
rect 109268 -972 109380 468
rect 110464 -972 110576 468
rect 111568 -972 111680 468
rect 112764 -972 112876 468
rect 113960 -972 114072 468
rect 115156 -972 115268 468
rect 116352 -972 116464 468
rect 117548 -972 117660 468
rect 118744 -972 118856 468
rect 119848 -972 119960 468
rect 121044 -972 121156 468
rect 122240 -972 122352 468
rect 123436 -972 123548 468
rect 124632 -972 124744 468
rect 125828 -972 125940 468
rect 126932 -972 127044 468
rect 128128 -972 128240 468
rect 129324 -972 129436 468
rect 130520 -972 130632 468
rect 131716 -972 131828 468
rect 132912 -972 133024 468
rect 134108 -972 134220 468
rect 135212 -972 135324 468
rect 136408 -972 136520 468
rect 137604 -972 137716 468
rect 138800 -972 138912 468
rect 139996 -972 140108 468
rect 141192 -972 141304 468
rect 142388 -972 142500 468
rect 143492 -972 143604 468
rect 144688 -972 144800 468
rect 145884 -972 145996 468
rect 147080 -972 147192 468
rect 148276 -972 148388 468
rect 149472 -972 149584 468
rect 150576 -972 150688 468
rect 151772 -972 151884 468
rect 152968 -972 153080 468
rect 154164 -972 154276 468
rect 155360 -972 155472 468
rect 156556 -972 156668 468
rect 157752 -972 157864 468
rect 158856 -972 158968 468
rect 160052 -972 160164 468
rect 161248 -972 161360 468
rect 162444 -972 162556 468
rect 163640 -972 163752 468
rect 164836 -972 164948 468
rect 166032 -972 166144 468
rect 167136 -972 167248 468
rect 168332 -972 168444 468
rect 169528 -972 169640 468
rect 170724 -972 170836 468
rect 171920 -972 172032 468
rect 173116 -972 173228 468
rect 174220 -972 174332 468
rect 175416 -972 175528 468
rect 176612 -972 176724 468
rect 177808 -972 177920 468
rect 179004 -972 179116 468
rect 180200 -972 180312 468
rect 181396 -972 181508 468
rect 182500 -972 182612 468
rect 183696 -972 183808 468
rect 184892 -972 185004 468
rect 186088 -972 186200 468
rect 187284 -972 187396 468
rect 188480 -972 188592 468
rect 189676 -972 189788 468
rect 190780 -972 190892 468
rect 191976 -972 192088 468
rect 193172 -972 193284 468
rect 194368 -972 194480 468
rect 195564 -972 195676 468
rect 196760 -972 196872 468
rect 197864 -972 197976 468
rect 199060 -972 199172 468
rect 200256 -972 200368 468
rect 201452 -972 201564 468
rect 202648 -972 202760 468
rect 203844 -972 203956 468
rect 205040 -972 205152 468
rect 206144 -972 206256 468
rect 207340 -972 207452 468
rect 208536 -972 208648 468
rect 209732 -972 209844 468
rect 210928 -972 211040 468
rect 212124 -972 212236 468
rect 213320 -972 213432 468
rect 214424 -972 214536 468
rect 215620 -972 215732 468
rect 216816 -972 216928 468
rect 218012 -972 218124 468
rect 219208 -972 219320 468
rect 220404 -972 220516 468
rect 221508 -972 221620 468
rect 222704 -972 222816 468
rect 223900 -972 224012 468
rect 225096 -972 225208 468
rect 226292 -972 226404 468
rect 227488 -972 227600 468
rect 228684 -972 228796 468
rect 229788 -972 229900 468
rect 230984 -972 231096 468
rect 232180 -972 232292 468
rect 233376 -972 233488 468
rect 234572 -972 234684 468
rect 235768 -972 235880 468
rect 236964 -972 237076 468
rect 238068 -972 238180 468
rect 239264 -972 239376 468
rect 240460 -972 240572 468
rect 241656 -972 241768 468
rect 242852 -972 242964 468
rect 244048 -972 244160 468
rect 245152 -972 245264 468
rect 246348 -972 246460 468
rect 247544 -972 247656 468
rect 248740 -972 248852 468
rect 249936 -972 250048 468
rect 251132 -972 251244 468
rect 252328 -972 252440 468
rect 253432 -972 253544 468
rect 254628 -972 254740 468
rect 255824 -972 255936 468
rect 257020 -972 257132 468
rect 258216 -972 258328 468
rect 259412 -972 259524 468
rect 260608 -972 260720 468
rect 261712 -972 261824 468
rect 262908 -972 263020 468
rect 264104 -972 264216 468
rect 265300 -972 265412 468
rect 266496 -972 266608 468
rect 267692 -972 267804 468
rect 268796 -972 268908 468
rect 269992 -972 270104 468
rect 271188 -972 271300 468
rect 272384 -972 272496 468
rect 273580 -972 273692 468
rect 274776 -972 274888 468
rect 275972 -972 276084 468
rect 277076 -972 277188 468
rect 278272 -972 278384 468
rect 279468 -972 279580 468
rect 280664 -972 280776 468
rect 281860 -972 281972 468
rect 283056 -972 283168 468
rect 284252 -972 284364 468
rect 285356 -972 285468 468
rect 286552 -972 286664 468
rect 287748 -972 287860 468
rect 288944 -972 289056 468
rect 290140 -972 290252 468
rect 291336 -972 291448 468
rect 292532 -972 292644 468
rect 293636 -972 293748 468
rect 294832 -972 294944 468
rect 296028 -972 296140 468
rect 297224 -972 297336 468
rect 298420 -972 298532 468
rect 299616 -972 299728 468
rect 300720 -972 300832 468
rect 301916 -972 302028 468
rect 303112 -972 303224 468
rect 304308 -972 304420 468
rect 305504 -972 305616 468
rect 306700 -972 306812 468
rect 307896 -972 308008 468
rect 309000 -972 309112 468
rect 310196 -972 310308 468
rect 311392 -972 311504 468
rect 312588 -972 312700 468
rect 313784 -972 313896 468
rect 314980 -972 315092 468
rect 316176 -972 316288 468
rect 317280 -972 317392 468
rect 318476 -972 318588 468
rect 319672 -972 319784 468
rect 320868 -972 320980 468
rect 322064 -972 322176 468
rect 323260 -972 323372 468
rect 324364 -972 324476 468
rect 325560 -972 325672 468
rect 326756 -972 326868 468
rect 327952 -972 328064 468
rect 329148 -972 329260 468
rect 330344 -972 330456 468
rect 331540 -972 331652 468
rect 332644 -972 332756 468
rect 333840 -972 333952 468
rect 335036 -972 335148 468
rect 336232 -972 336344 468
rect 337428 -972 337540 468
rect 338624 -972 338736 468
rect 339820 -972 339932 468
rect 340924 -972 341036 468
rect 342120 -972 342232 468
rect 343316 -972 343428 468
rect 344512 -972 344624 468
rect 345708 -972 345820 468
rect 346904 -972 347016 468
rect 348008 -972 348120 468
rect 349204 -972 349316 468
rect 350400 -972 350512 468
rect 351596 -972 351708 468
rect 352792 -972 352904 468
rect 353988 -972 354100 468
rect 355184 -972 355296 468
rect 356288 -972 356400 468
rect 357484 -972 357596 468
rect 358680 -972 358792 468
rect 359876 -972 359988 468
rect 361072 -972 361184 468
rect 362268 -972 362380 468
rect 363464 -972 363576 468
rect 364568 -972 364680 468
rect 365764 -972 365876 468
rect 366960 -972 367072 468
rect 368156 -972 368268 468
rect 369352 -972 369464 468
rect 370548 -972 370660 468
rect 371652 -972 371764 468
rect 372848 -972 372960 468
rect 374044 -972 374156 468
rect 375240 -972 375352 468
rect 376436 -972 376548 468
rect 377632 -972 377744 468
rect 378828 -972 378940 468
rect 379932 -972 380044 468
rect 381128 -972 381240 468
rect 382324 -972 382436 468
rect 383520 -972 383632 468
rect 384716 -972 384828 468
rect 385912 -972 386024 468
rect 387108 -972 387220 468
rect 388212 -972 388324 468
rect 389408 -972 389520 468
rect 390604 -972 390716 468
rect 391800 -972 391912 468
rect 392996 -972 393108 468
rect 394192 -972 394304 468
rect 395296 -972 395408 468
rect 396492 -972 396604 468
rect 397688 -972 397800 468
rect 398884 -972 398996 468
rect 400080 -972 400192 468
rect 401276 -972 401388 468
rect 402472 -972 402584 468
rect 403576 -972 403688 468
rect 404772 -972 404884 468
rect 405968 -972 406080 468
rect 407164 -972 407276 468
rect 408360 -972 408472 468
rect 409556 -972 409668 468
rect 410752 -972 410864 468
rect 411856 -972 411968 468
rect 413052 -972 413164 468
rect 414248 -972 414360 468
rect 415444 -972 415556 468
rect 416640 -972 416752 468
rect 417836 -972 417948 468
rect 418940 -972 419052 468
rect 420136 -972 420248 468
rect 421332 -972 421444 468
rect 422528 -972 422640 468
rect 423724 -972 423836 468
rect 424920 -972 425032 468
rect 426116 -972 426228 468
rect 427220 -972 427332 468
rect 428416 -972 428528 468
rect 429612 -972 429724 468
rect 430808 -972 430920 468
rect 432004 -972 432116 468
rect 433200 -972 433312 468
rect 434396 -972 434508 468
rect 435500 -972 435612 468
rect 436696 -972 436808 468
rect 437892 -972 438004 468
rect 439088 -972 439200 468
rect 440284 -972 440396 468
rect 441480 -972 441592 468
rect 442584 -972 442696 468
rect 443780 -972 443892 468
rect 444976 -972 445088 468
rect 446172 -972 446284 468
rect 447368 -972 447480 468
rect 448564 -972 448676 468
rect 449760 -972 449872 468
rect 450864 -972 450976 468
rect 452060 -972 452172 468
rect 453256 -972 453368 468
rect 454452 -972 454564 468
rect 455648 -972 455760 468
rect 456844 -972 456956 468
rect 458040 -972 458152 468
rect 459144 -972 459256 468
rect 460340 -972 460452 468
rect 461536 -972 461648 468
rect 462732 -972 462844 468
rect 463928 -972 464040 468
rect 465124 -972 465236 468
rect 466228 -972 466340 468
rect 467424 -972 467536 468
rect 468620 -972 468732 468
rect 469816 -972 469928 468
rect 471012 -972 471124 468
rect 472208 -972 472320 468
rect 473404 -972 473516 468
rect 474508 -972 474620 468
rect 475704 -972 475816 468
rect 476900 -972 477012 468
rect 478096 -972 478208 468
rect 479292 -972 479404 468
rect 480488 -972 480600 468
rect 481684 -972 481796 468
rect 482788 -972 482900 468
rect 483984 -972 484096 468
rect 485180 -972 485292 468
rect 486376 -972 486488 468
rect 487572 -972 487684 468
rect 488768 -972 488880 468
rect 489872 -972 489984 468
rect 491068 -972 491180 468
rect 492264 -972 492376 468
rect 493460 -972 493572 468
rect 494656 -972 494768 468
rect 495852 -972 495964 468
rect 497048 -972 497160 468
rect 498152 -972 498264 468
rect 499348 -972 499460 468
rect 500544 -972 500656 468
rect 501740 -972 501852 468
rect 502936 -972 503048 468
rect 504132 -972 504244 468
rect 505328 -972 505440 468
rect 506432 -972 506544 468
rect 507628 -972 507740 468
rect 508824 -972 508936 468
rect 510020 -972 510132 468
rect 511216 -972 511328 468
rect 512412 -972 512524 468
rect 513516 -972 513628 468
rect 514712 -972 514824 468
rect 515908 -972 516020 468
rect 517104 -972 517216 468
rect 518300 -972 518412 468
rect 519496 -972 519608 468
rect 520692 -972 520804 468
rect 521796 -972 521908 468
rect 522992 -972 523104 468
rect 524188 -972 524300 468
rect 525384 -972 525496 468
rect 526580 -972 526692 468
rect 527776 -972 527888 468
rect 528972 -972 529084 468
rect 530076 -972 530188 468
rect 531272 -972 531384 468
rect 532468 -972 532580 468
rect 533664 -972 533776 468
rect 534860 -972 534972 468
rect 536056 -972 536168 468
rect 537160 -972 537272 468
rect 538356 -972 538468 468
rect 539552 -972 539664 468
rect 540748 -972 540860 468
rect 541944 -972 542056 468
rect 543140 -972 543252 468
rect 544336 -972 544448 468
rect 545440 -972 545552 468
rect 546636 -972 546748 468
rect 547832 -972 547944 468
rect 549028 -972 549140 468
rect 550224 -972 550336 468
rect 551420 -972 551532 468
rect 552616 -972 552728 468
rect 553720 -972 553832 468
rect 554916 -972 555028 468
rect 556112 -972 556224 468
rect 557308 -972 557420 468
rect 558504 -972 558616 468
rect 559700 -972 559812 468
rect 560804 -972 560916 468
rect 562000 -972 562112 468
rect 563196 -972 563308 468
rect 564392 -972 564504 468
rect 565588 -972 565700 468
rect 566784 -972 566896 468
rect 567980 -972 568092 468
rect 569084 -972 569196 468
rect 570280 -972 570392 468
rect 571476 -972 571588 468
rect 572672 -972 572784 468
rect 573868 -972 573980 468
rect 575064 -972 575176 468
rect 576260 -972 576372 468
rect 577364 -972 577476 468
rect 578560 -972 578672 468
rect 579756 -972 579868 468
rect 580952 -972 581064 468
rect 582148 -972 582260 468
rect 583344 -972 583456 468
<< via2 >>
rect 351424 626932 351850 628628
rect 371240 644684 372084 644874
rect 372762 644690 373386 644868
rect 370660 641480 371192 641666
rect 373272 641496 373888 641664
rect 371028 636912 371560 637098
rect 373040 636928 373656 637096
rect 371548 624430 371696 625304
rect 372000 624060 372174 624632
rect 372782 624080 372956 624652
rect 371568 622312 371742 622884
<< metal3 >>
rect -978 698976 462 699216
rect 583502 698840 584942 699080
rect -978 689592 372570 689832
rect -978 680208 462 680448
rect -978 670824 462 671064
rect -978 661440 462 661680
rect -978 652056 462 652296
rect 371198 644874 372122 644900
rect 371198 644684 371240 644874
rect 372084 644870 372122 644874
rect 372084 644684 372126 644870
rect 371198 644650 372126 644684
rect 371200 644648 372126 644650
rect -978 642672 462 642912
rect 370616 641666 371248 641698
rect 370616 641574 370660 641666
rect 370522 641566 370660 641574
rect 351100 641506 370660 641566
rect -978 633288 462 633528
rect 351100 624480 351160 641506
rect 370488 641505 370660 641506
rect 370616 641480 370660 641505
rect 371192 641480 371248 641666
rect 370616 641454 371248 641480
rect 371940 640150 372000 644648
rect 352265 640090 372000 640150
rect 351354 628628 351968 628750
rect 351354 626932 351424 628628
rect 351850 626932 351968 628628
rect 351354 626848 351968 626932
rect 350044 624420 351160 624480
rect -978 623904 462 624144
rect 352265 624115 352325 640090
rect 370984 637098 371616 637130
rect 370984 637006 371028 637098
rect 350044 624055 352325 624115
rect 352582 636937 371028 637006
rect 352582 623398 352651 636937
rect 370984 636912 371028 636937
rect 371560 636912 371616 637098
rect 370984 636886 371616 636912
rect 371484 625304 371740 625348
rect 371484 624472 371548 625304
rect 364168 624430 371548 624472
rect 371696 624430 371740 625304
rect 364168 624412 371740 624430
rect 371484 624378 371740 624412
rect 371972 624632 372212 624672
rect 371972 624107 372000 624632
rect 364168 624060 372000 624107
rect 372174 624060 372212 624632
rect 364168 624047 372212 624060
rect 371972 624002 372212 624047
rect 350044 623329 352651 623398
rect 372330 623390 372570 689592
rect 583502 688912 584942 689152
rect 583502 678984 584942 679224
rect 583502 669056 584942 669296
rect 583502 659128 584942 659368
rect 583502 649200 584942 649440
rect 372714 644868 400212 644894
rect 372714 644690 372762 644868
rect 373386 644690 400212 644868
rect 372714 644654 400212 644690
rect 373226 641664 396442 641718
rect 373226 641496 373272 641664
rect 373888 641496 396442 641664
rect 373226 641478 396442 641496
rect 373226 641452 374210 641478
rect 372986 637096 389758 637124
rect 372986 636928 373040 637096
rect 373656 636928 389758 637096
rect 372986 636884 389758 636928
rect 372754 624652 372994 624692
rect 372754 624080 372782 624652
rect 372956 624184 372994 624652
rect 372956 624080 377900 624184
rect 372754 624052 377900 624080
rect 372754 624022 372994 624052
rect 364168 623322 372570 623390
rect 364168 623321 372558 623322
rect 371540 622884 371780 622924
rect 371540 622312 371568 622884
rect 371742 622312 371780 622884
rect -978 614520 462 614760
rect -978 605136 462 605376
rect -978 595752 462 595992
rect -978 586368 462 586608
rect 371540 577224 371780 622312
rect -978 576984 371780 577224
rect -978 567600 462 567840
rect -978 558216 462 558456
rect -978 548832 462 549072
rect -978 539448 462 539688
rect -978 530064 462 530304
rect 377660 520920 377900 624052
rect -978 520680 377900 520920
rect -978 511296 462 511536
rect -978 501912 462 502152
rect -978 492528 462 492768
rect -978 483144 462 483384
rect -978 473760 462 474000
rect -978 464376 462 464616
rect 389518 461080 389758 636884
rect 396202 560224 396442 641478
rect 399972 619656 400212 644654
rect 583502 639272 584942 639512
rect 583502 629344 584942 629584
rect 399972 619416 584942 619656
rect 583502 609488 584942 609728
rect 583502 599696 584942 599936
rect 583502 589768 584942 590008
rect 583502 579840 584942 580080
rect 583502 569912 584942 570152
rect 396202 559984 584942 560224
rect 583502 550056 584942 550296
rect 583502 540128 584942 540368
rect 583502 530200 584942 530440
rect 583502 520272 584942 520512
rect 583502 510344 584942 510584
rect 583502 500552 584942 500792
rect 583502 490624 584942 490864
rect 583502 480696 584942 480936
rect 583502 470768 584942 471008
rect 389518 460840 584942 461080
rect -978 454992 462 455232
rect 583502 450912 584942 451152
rect -978 445608 462 445848
rect 583502 440984 584942 441224
rect -978 436224 462 436464
rect 583502 431056 584942 431296
rect -978 426840 462 427080
rect 583502 421128 584942 421368
rect -978 417456 462 417696
rect 583502 411200 584942 411440
rect -978 408072 462 408312
rect 583502 401408 584942 401648
rect -978 398688 462 398928
rect 583502 391480 584942 391720
rect -978 389304 462 389544
rect 583502 381552 584942 381792
rect -978 379920 462 380160
rect 583502 371624 584942 371864
rect -978 370536 462 370776
rect 583502 361696 584942 361936
rect -978 361152 462 361392
rect -978 351768 462 352008
rect 583502 351768 584942 352008
rect -978 342384 462 342624
rect 583502 341840 584942 342080
rect -978 333000 462 333240
rect 583502 331912 584942 332152
rect -978 323616 462 323856
rect 583502 321984 584942 322224
rect -978 314232 462 314472
rect 583502 312056 584942 312296
rect -978 304848 462 305088
rect 583502 302264 584942 302504
rect -978 295464 462 295704
rect 583502 292336 584942 292576
rect -978 286080 462 286320
rect 583502 282408 584942 282648
rect -978 276696 462 276936
rect 583502 272480 584942 272720
rect -978 267312 462 267552
rect 583502 262552 584942 262792
rect -978 257928 462 258168
rect 583502 252624 584942 252864
rect -978 248544 462 248784
rect 583502 242696 584942 242936
rect -978 239160 462 239400
rect 583502 232768 584942 233008
rect -978 229776 462 230016
rect 583502 222840 584942 223080
rect -978 220392 462 220632
rect 583502 212912 584942 213152
rect -978 211008 462 211248
rect 583502 203120 584942 203360
rect -978 201624 462 201864
rect 583502 193192 584942 193432
rect -978 192240 462 192480
rect 583502 183264 584942 183504
rect -978 182856 462 183096
rect -978 173472 462 173712
rect 583502 173336 584942 173576
rect -978 164088 462 164328
rect 583502 163408 584942 163648
rect -978 154704 462 154944
rect 583502 153480 584942 153720
rect -978 145320 462 145560
rect 583502 143552 584942 143792
rect -978 135936 462 136176
rect 583502 133624 584942 133864
rect -978 126552 462 126792
rect 583502 123696 584942 123936
rect -978 117168 462 117408
rect 583502 113768 584942 114008
rect -978 107784 462 108024
rect 583502 103976 584942 104216
rect -978 98400 462 98640
rect 583502 94048 584942 94288
rect -978 89016 462 89256
rect 583502 84120 584942 84360
rect -978 79632 462 79872
rect 583502 74192 584942 74432
rect -978 70248 462 70488
rect 583502 64264 584942 64504
rect -978 60864 462 61104
rect 583502 54336 584942 54576
rect -978 51480 462 51720
rect 583502 44408 584942 44648
rect -978 42096 462 42336
rect 583502 34480 584942 34720
rect -978 32712 462 32952
rect 583502 24552 584942 24792
rect -978 23328 462 23568
rect 583502 14624 584942 14864
rect -978 13944 462 14184
rect 583502 4832 584942 5072
rect -978 4560 462 4800
<< via3 >>
rect 351424 626932 351850 628628
<< metal4 >>
rect -8594 711406 -7994 711428
rect -8594 711170 -8412 711406
rect -8176 711170 -7994 711406
rect -8594 711086 -7994 711170
rect -8594 710850 -8412 711086
rect -8176 710850 -7994 711086
rect -8594 -6938 -7994 710850
rect 591882 711406 592482 711428
rect 591882 711170 592064 711406
rect 592300 711170 592482 711406
rect 591882 711086 592482 711170
rect 591882 710850 592064 711086
rect 592300 710850 592482 711086
rect -7654 710466 -7054 710488
rect -7654 710230 -7472 710466
rect -7236 710230 -7054 710466
rect -7654 710146 -7054 710230
rect -7654 709910 -7472 710146
rect -7236 709910 -7054 710146
rect -7654 -5998 -7054 709910
rect 590942 710466 591542 710488
rect 590942 710230 591124 710466
rect 591360 710230 591542 710466
rect 590942 710146 591542 710230
rect 590942 709910 591124 710146
rect 591360 709910 591542 710146
rect -6714 709526 -6114 709548
rect -6714 709290 -6532 709526
rect -6296 709290 -6114 709526
rect -6714 709206 -6114 709290
rect -6714 708970 -6532 709206
rect -6296 708970 -6114 709206
rect -6714 -5058 -6114 708970
rect 343100 709500 344038 709618
rect 343100 708996 343160 709500
rect 343966 708996 344038 709500
rect -5774 708586 -5174 708608
rect -5774 708350 -5592 708586
rect -5356 708350 -5174 708586
rect -5774 708266 -5174 708350
rect -5774 708030 -5592 708266
rect -5356 708030 -5174 708266
rect -5774 -4118 -5174 708030
rect -4834 707646 -4234 707668
rect -4834 707410 -4652 707646
rect -4416 707410 -4234 707646
rect -4834 707326 -4234 707410
rect -4834 707090 -4652 707326
rect -4416 707090 -4234 707326
rect -4834 -3178 -4234 707090
rect -3894 706706 -3294 706728
rect -3894 706470 -3712 706706
rect -3476 706470 -3294 706706
rect -3894 706386 -3294 706470
rect -3894 706150 -3712 706386
rect -3476 706150 -3294 706386
rect -3894 -2238 -3294 706150
rect -2954 705766 -2354 705788
rect -2954 705530 -2772 705766
rect -2536 705530 -2354 705766
rect -2954 705446 -2354 705530
rect -2954 705210 -2772 705446
rect -2536 705210 -2354 705446
rect -2954 -1298 -2354 705210
rect -2014 704826 -1414 704848
rect -2014 704590 -1832 704826
rect -1596 704590 -1414 704826
rect -2014 704506 -1414 704590
rect -2014 704270 -1832 704506
rect -1596 704270 -1414 704506
rect -2014 -358 -1414 704270
rect 343100 698930 344038 708996
rect 357218 709494 358156 709588
rect 357218 708990 357280 709494
rect 358086 708990 358156 709494
rect 351430 708596 351846 708622
rect 351138 708524 352174 708596
rect 351138 708076 351240 708524
rect 352044 708076 352174 708524
rect 351138 708018 352174 708076
rect 350523 704806 350852 704880
rect 350523 704288 350554 704806
rect 350816 704288 350852 704806
rect 350523 624855 350852 704288
rect 351430 630020 351846 708018
rect 357218 699046 358156 708990
rect 590002 709526 590602 709548
rect 590002 709290 590184 709526
rect 590420 709290 590602 709526
rect 590002 709206 590602 709290
rect 590002 708970 590184 709206
rect 590420 708970 590602 709206
rect 589062 708586 589662 708608
rect 589062 708350 589244 708586
rect 589480 708350 589662 708586
rect 589062 708266 589662 708350
rect 589062 708030 589244 708266
rect 589480 708030 589662 708266
rect 588122 707646 588722 707668
rect 588122 707410 588304 707646
rect 588540 707410 588722 707646
rect 588122 707326 588722 707410
rect 588122 707090 588304 707326
rect 588540 707090 588722 707326
rect 587182 706706 587782 706728
rect 587182 706470 587364 706706
rect 587600 706470 587782 706706
rect 587182 706386 587782 706470
rect 587182 706150 587364 706386
rect 587600 706150 587782 706386
rect 586242 705766 586842 705788
rect 586242 705530 586424 705766
rect 586660 705530 586842 705766
rect 586242 705446 586842 705530
rect 586242 705210 586424 705446
rect 586660 705210 586842 705446
rect 365282 704818 365616 704864
rect 365282 704272 365304 704818
rect 365596 704272 365616 704818
rect 351432 628750 351844 630020
rect 351354 628628 351968 628750
rect 351354 626932 351424 628628
rect 351850 626932 351968 628628
rect 365282 628604 365616 704272
rect 585302 704826 585902 704848
rect 585302 704590 585484 704826
rect 585720 704590 585902 704826
rect 585302 704506 585902 704590
rect 585302 704270 585484 704506
rect 585720 704270 585902 704506
rect 351354 626848 351968 626932
rect 349828 624526 350858 624855
rect 365285 624847 365614 628604
rect 364046 624518 365614 624847
rect -2014 -594 -1832 -358
rect -1596 -594 -1414 -358
rect -2014 -678 -1414 -594
rect -2014 -914 -1832 -678
rect -1596 -914 -1414 -678
rect -2014 -936 -1414 -914
rect 585302 -358 585902 704270
rect 585302 -594 585484 -358
rect 585720 -594 585902 -358
rect 585302 -678 585902 -594
rect 585302 -914 585484 -678
rect 585720 -914 585902 -678
rect 585302 -936 585902 -914
rect -2954 -1534 -2772 -1298
rect -2536 -1534 -2354 -1298
rect -2954 -1618 -2354 -1534
rect -2954 -1854 -2772 -1618
rect -2536 -1854 -2354 -1618
rect -2954 -1876 -2354 -1854
rect 586242 -1298 586842 705210
rect 586242 -1534 586424 -1298
rect 586660 -1534 586842 -1298
rect 586242 -1618 586842 -1534
rect 586242 -1854 586424 -1618
rect 586660 -1854 586842 -1618
rect 586242 -1876 586842 -1854
rect -3894 -2474 -3712 -2238
rect -3476 -2474 -3294 -2238
rect -3894 -2558 -3294 -2474
rect -3894 -2794 -3712 -2558
rect -3476 -2794 -3294 -2558
rect -3894 -2816 -3294 -2794
rect 587182 -2238 587782 706150
rect 587182 -2474 587364 -2238
rect 587600 -2474 587782 -2238
rect 587182 -2558 587782 -2474
rect 587182 -2794 587364 -2558
rect 587600 -2794 587782 -2558
rect 587182 -2816 587782 -2794
rect -4834 -3414 -4652 -3178
rect -4416 -3414 -4234 -3178
rect -4834 -3498 -4234 -3414
rect -4834 -3734 -4652 -3498
rect -4416 -3734 -4234 -3498
rect -4834 -3756 -4234 -3734
rect 588122 -3178 588722 707090
rect 588122 -3414 588304 -3178
rect 588540 -3414 588722 -3178
rect 588122 -3498 588722 -3414
rect 588122 -3734 588304 -3498
rect 588540 -3734 588722 -3498
rect 588122 -3756 588722 -3734
rect -5774 -4354 -5592 -4118
rect -5356 -4354 -5174 -4118
rect -5774 -4438 -5174 -4354
rect -5774 -4674 -5592 -4438
rect -5356 -4674 -5174 -4438
rect -5774 -4696 -5174 -4674
rect 589062 -4118 589662 708030
rect 589062 -4354 589244 -4118
rect 589480 -4354 589662 -4118
rect 589062 -4438 589662 -4354
rect 589062 -4674 589244 -4438
rect 589480 -4674 589662 -4438
rect 589062 -4696 589662 -4674
rect -6714 -5294 -6532 -5058
rect -6296 -5294 -6114 -5058
rect -6714 -5378 -6114 -5294
rect -6714 -5614 -6532 -5378
rect -6296 -5614 -6114 -5378
rect -6714 -5636 -6114 -5614
rect 590002 -5058 590602 708970
rect 590002 -5294 590184 -5058
rect 590420 -5294 590602 -5058
rect 590002 -5378 590602 -5294
rect 590002 -5614 590184 -5378
rect 590420 -5614 590602 -5378
rect 590002 -5636 590602 -5614
rect -7654 -6234 -7472 -5998
rect -7236 -6234 -7054 -5998
rect -7654 -6318 -7054 -6234
rect -7654 -6554 -7472 -6318
rect -7236 -6554 -7054 -6318
rect -7654 -6576 -7054 -6554
rect 590942 -5998 591542 709910
rect 590942 -6234 591124 -5998
rect 591360 -6234 591542 -5998
rect 590942 -6318 591542 -6234
rect 590942 -6554 591124 -6318
rect 591360 -6554 591542 -6318
rect 590942 -6576 591542 -6554
rect -8594 -7174 -8412 -6938
rect -8176 -7174 -7994 -6938
rect -8594 -7258 -7994 -7174
rect -8594 -7494 -8412 -7258
rect -8176 -7494 -7994 -7258
rect -8594 -7516 -7994 -7494
rect 591882 -6938 592482 710850
rect 591882 -7174 592064 -6938
rect 592300 -7174 592482 -6938
rect 591882 -7258 592482 -7174
rect 591882 -7494 592064 -7258
rect 592300 -7494 592482 -7258
rect 591882 -7516 592482 -7494
<< via4 >>
rect -8412 711170 -8176 711406
rect -8412 710850 -8176 711086
rect 592064 711170 592300 711406
rect 592064 710850 592300 711086
rect -7472 710230 -7236 710466
rect -7472 709910 -7236 710146
rect 591124 710230 591360 710466
rect 591124 709910 591360 710146
rect -6532 709290 -6296 709526
rect -6532 708970 -6296 709206
rect 343160 708996 343966 709500
rect -5592 708350 -5356 708586
rect -5592 708030 -5356 708266
rect -4652 707410 -4416 707646
rect -4652 707090 -4416 707326
rect -3712 706470 -3476 706706
rect -3712 706150 -3476 706386
rect -2772 705530 -2536 705766
rect -2772 705210 -2536 705446
rect -1832 704590 -1596 704826
rect -1832 704270 -1596 704506
rect 357280 708990 358086 709494
rect 351240 708076 352044 708524
rect 350554 704288 350816 704806
rect 590184 709290 590420 709526
rect 590184 708970 590420 709206
rect 589244 708350 589480 708586
rect 589244 708030 589480 708266
rect 588304 707410 588540 707646
rect 588304 707090 588540 707326
rect 587364 706470 587600 706706
rect 587364 706150 587600 706386
rect 586424 705530 586660 705766
rect 586424 705210 586660 705446
rect 365304 704272 365596 704818
rect 585484 704590 585720 704826
rect 585484 704270 585720 704506
rect -1832 -594 -1596 -358
rect -1832 -914 -1596 -678
rect 585484 -594 585720 -358
rect 585484 -914 585720 -678
rect -2772 -1534 -2536 -1298
rect -2772 -1854 -2536 -1618
rect 586424 -1534 586660 -1298
rect 586424 -1854 586660 -1618
rect -3712 -2474 -3476 -2238
rect -3712 -2794 -3476 -2558
rect 587364 -2474 587600 -2238
rect 587364 -2794 587600 -2558
rect -4652 -3414 -4416 -3178
rect -4652 -3734 -4416 -3498
rect 588304 -3414 588540 -3178
rect 588304 -3734 588540 -3498
rect -5592 -4354 -5356 -4118
rect -5592 -4674 -5356 -4438
rect 589244 -4354 589480 -4118
rect 589244 -4674 589480 -4438
rect -6532 -5294 -6296 -5058
rect -6532 -5614 -6296 -5378
rect 590184 -5294 590420 -5058
rect 590184 -5614 590420 -5378
rect -7472 -6234 -7236 -5998
rect -7472 -6554 -7236 -6318
rect 591124 -6234 591360 -5998
rect 591124 -6554 591360 -6318
rect -8412 -7174 -8176 -6938
rect -8412 -7494 -8176 -7258
rect 592064 -7174 592300 -6938
rect 592064 -7494 592300 -7258
<< metal5 >>
rect -8594 711428 -7994 711430
rect 591882 711428 592482 711430
rect -8594 711406 592482 711428
rect -8594 711170 -8412 711406
rect -8176 711170 592064 711406
rect 592300 711170 592482 711406
rect -8594 711086 592482 711170
rect -8594 710850 -8412 711086
rect -8176 710850 592064 711086
rect 592300 710850 592482 711086
rect -8594 710828 592482 710850
rect -8594 710826 -7994 710828
rect 591882 710826 592482 710828
rect -7654 710488 -7054 710490
rect 590942 710488 591542 710490
rect -7654 710466 591542 710488
rect -7654 710230 -7472 710466
rect -7236 710230 591124 710466
rect 591360 710230 591542 710466
rect -7654 710146 591542 710230
rect -7654 709910 -7472 710146
rect -7236 709910 591124 710146
rect 591360 709910 591542 710146
rect -7654 709888 591542 709910
rect -7654 709886 -7054 709888
rect 590942 709886 591542 709888
rect -6714 709548 -6114 709550
rect 590002 709548 590602 709550
rect -6714 709526 590602 709548
rect -6714 709290 -6532 709526
rect -6296 709500 590184 709526
rect -6296 709290 343160 709500
rect -6714 709206 343160 709290
rect -6714 708970 -6532 709206
rect -6296 708996 343160 709206
rect 343966 709494 590184 709500
rect 343966 708996 357280 709494
rect -6296 708990 357280 708996
rect 358086 709290 590184 709494
rect 590420 709290 590602 709526
rect 358086 709206 590602 709290
rect 358086 708990 590184 709206
rect -6296 708970 590184 708990
rect 590420 708970 590602 709206
rect -6714 708948 590602 708970
rect -6714 708946 -6114 708948
rect 590002 708946 590602 708948
rect -5774 708608 -5174 708610
rect 589062 708608 589662 708610
rect -5774 708586 589662 708608
rect -5774 708350 -5592 708586
rect -5356 708524 589244 708586
rect -5356 708350 351240 708524
rect -5774 708266 351240 708350
rect -5774 708030 -5592 708266
rect -5356 708076 351240 708266
rect 352044 708350 589244 708524
rect 589480 708350 589662 708586
rect 352044 708266 589662 708350
rect 352044 708076 589244 708266
rect -5356 708030 589244 708076
rect 589480 708030 589662 708266
rect -5774 708008 589662 708030
rect -5774 708006 -5174 708008
rect 589062 708006 589662 708008
rect -4834 707668 -4234 707670
rect 588122 707668 588722 707670
rect -4834 707646 588722 707668
rect -4834 707410 -4652 707646
rect -4416 707410 588304 707646
rect 588540 707410 588722 707646
rect -4834 707326 588722 707410
rect -4834 707090 -4652 707326
rect -4416 707090 588304 707326
rect 588540 707090 588722 707326
rect -4834 707068 588722 707090
rect -4834 707066 -4234 707068
rect 588122 707066 588722 707068
rect -3894 706728 -3294 706730
rect 587182 706728 587782 706730
rect -3894 706706 587782 706728
rect -3894 706470 -3712 706706
rect -3476 706470 587364 706706
rect 587600 706470 587782 706706
rect -3894 706386 587782 706470
rect -3894 706150 -3712 706386
rect -3476 706150 587364 706386
rect 587600 706150 587782 706386
rect -3894 706128 587782 706150
rect -3894 706126 -3294 706128
rect 587182 706126 587782 706128
rect -2954 705788 -2354 705790
rect 586242 705788 586842 705790
rect -2954 705766 586842 705788
rect -2954 705530 -2772 705766
rect -2536 705530 586424 705766
rect 586660 705530 586842 705766
rect -2954 705446 586842 705530
rect -2954 705210 -2772 705446
rect -2536 705210 586424 705446
rect 586660 705210 586842 705446
rect -2954 705188 586842 705210
rect -2954 705186 -2354 705188
rect 586242 705186 586842 705188
rect -2014 704848 -1414 704850
rect 585302 704848 585902 704850
rect -2014 704826 585902 704848
rect -2014 704590 -1832 704826
rect -1596 704818 585484 704826
rect -1596 704806 365304 704818
rect -1596 704590 350554 704806
rect -2014 704506 350554 704590
rect -2014 704270 -1832 704506
rect -1596 704288 350554 704506
rect 350816 704288 365304 704806
rect -1596 704272 365304 704288
rect 365596 704590 585484 704818
rect 585720 704590 585902 704826
rect 365596 704506 585902 704590
rect 365596 704272 585484 704506
rect -1596 704270 585484 704272
rect 585720 704270 585902 704506
rect -2014 704248 585902 704270
rect -2014 704246 -1414 704248
rect 585302 704246 585902 704248
rect 343130 623776 344004 701299
rect 357252 623768 358152 702284
rect -2014 -336 -1414 -334
rect 585302 -336 585902 -334
rect -2014 -358 585902 -336
rect -2014 -594 -1832 -358
rect -1596 -594 585484 -358
rect 585720 -594 585902 -358
rect -2014 -678 585902 -594
rect -2014 -914 -1832 -678
rect -1596 -914 585484 -678
rect 585720 -914 585902 -678
rect -2014 -936 585902 -914
rect -2014 -938 -1414 -936
rect 585302 -938 585902 -936
rect -2954 -1276 -2354 -1274
rect 586242 -1276 586842 -1274
rect -2954 -1298 586842 -1276
rect -2954 -1534 -2772 -1298
rect -2536 -1534 586424 -1298
rect 586660 -1534 586842 -1298
rect -2954 -1618 586842 -1534
rect -2954 -1854 -2772 -1618
rect -2536 -1854 586424 -1618
rect 586660 -1854 586842 -1618
rect -2954 -1876 586842 -1854
rect -2954 -1878 -2354 -1876
rect 586242 -1878 586842 -1876
rect -3894 -2216 -3294 -2214
rect 587182 -2216 587782 -2214
rect -3894 -2238 587782 -2216
rect -3894 -2474 -3712 -2238
rect -3476 -2474 587364 -2238
rect 587600 -2474 587782 -2238
rect -3894 -2558 587782 -2474
rect -3894 -2794 -3712 -2558
rect -3476 -2794 587364 -2558
rect 587600 -2794 587782 -2558
rect -3894 -2816 587782 -2794
rect -3894 -2818 -3294 -2816
rect 587182 -2818 587782 -2816
rect -4834 -3156 -4234 -3154
rect 588122 -3156 588722 -3154
rect -4834 -3178 588722 -3156
rect -4834 -3414 -4652 -3178
rect -4416 -3414 588304 -3178
rect 588540 -3414 588722 -3178
rect -4834 -3498 588722 -3414
rect -4834 -3734 -4652 -3498
rect -4416 -3734 588304 -3498
rect 588540 -3734 588722 -3498
rect -4834 -3756 588722 -3734
rect -4834 -3758 -4234 -3756
rect 588122 -3758 588722 -3756
rect -5774 -4096 -5174 -4094
rect 589062 -4096 589662 -4094
rect -5774 -4118 589662 -4096
rect -5774 -4354 -5592 -4118
rect -5356 -4354 589244 -4118
rect 589480 -4354 589662 -4118
rect -5774 -4438 589662 -4354
rect -5774 -4674 -5592 -4438
rect -5356 -4674 589244 -4438
rect 589480 -4674 589662 -4438
rect -5774 -4696 589662 -4674
rect -5774 -4698 -5174 -4696
rect 589062 -4698 589662 -4696
rect -6714 -5036 -6114 -5034
rect 590002 -5036 590602 -5034
rect -6714 -5058 590602 -5036
rect -6714 -5294 -6532 -5058
rect -6296 -5294 590184 -5058
rect 590420 -5294 590602 -5058
rect -6714 -5378 590602 -5294
rect -6714 -5614 -6532 -5378
rect -6296 -5614 590184 -5378
rect 590420 -5614 590602 -5378
rect -6714 -5636 590602 -5614
rect -6714 -5638 -6114 -5636
rect 590002 -5638 590602 -5636
rect -7654 -5976 -7054 -5974
rect 590942 -5976 591542 -5974
rect -7654 -5998 591542 -5976
rect -7654 -6234 -7472 -5998
rect -7236 -6234 591124 -5998
rect 591360 -6234 591542 -5998
rect -7654 -6318 591542 -6234
rect -7654 -6554 -7472 -6318
rect -7236 -6554 591124 -6318
rect 591360 -6554 591542 -6318
rect -7654 -6576 591542 -6554
rect -7654 -6578 -7054 -6576
rect 590942 -6578 591542 -6576
rect -8594 -6916 -7994 -6914
rect 591882 -6916 592482 -6914
rect -8594 -6938 592482 -6916
rect -8594 -7174 -8412 -6938
rect -8176 -7174 592064 -6938
rect 592300 -7174 592482 -6938
rect -8594 -7258 592482 -7174
rect -8594 -7494 -8412 -7258
rect -8176 -7494 592064 -7258
rect 592300 -7494 592482 -7258
rect -8594 -7516 592482 -7494
rect -8594 -7518 -7994 -7516
rect 591882 -7518 592482 -7516
use user_analog_proj_example  user_analog_proj_example_0
timestamp 1619730755
transform 1 0 338772 0 1 616578
box -26 -22 25476 8324
<< labels >>
rlabel metal3 s 583502 282408 584942 282648 6 gpio_analog[0]
port 0 nsew signal bidirectional
rlabel metal3 s -978 558216 462 558456 4 gpio_analog[10]
port 1 nsew signal bidirectional
rlabel metal3 s -978 501912 462 502152 4 gpio_analog[11]
port 2 nsew signal bidirectional
rlabel metal3 s -978 445608 462 445848 4 gpio_analog[12]
port 3 nsew signal bidirectional
rlabel metal3 s -978 389304 462 389544 4 gpio_analog[13]
port 4 nsew signal bidirectional
rlabel metal3 s -978 333000 462 333240 4 gpio_analog[14]
port 5 nsew signal bidirectional
rlabel metal3 s -978 276696 462 276936 4 gpio_analog[15]
port 6 nsew signal bidirectional
rlabel metal3 s -978 220392 462 220632 4 gpio_analog[16]
port 7 nsew signal bidirectional
rlabel metal3 s -978 164088 462 164328 4 gpio_analog[17]
port 8 nsew signal bidirectional
rlabel metal3 s 583502 341840 584942 342080 6 gpio_analog[1]
port 9 nsew signal bidirectional
rlabel metal3 s 583502 401408 584942 401648 6 gpio_analog[2]
port 10 nsew signal bidirectional
rlabel metal3 s 583502 460840 584942 461080 6 gpio_analog[3]
port 11 nsew signal bidirectional
rlabel metal3 s 583502 520272 584942 520512 6 gpio_analog[4]
port 12 nsew signal bidirectional
rlabel metal3 s 583502 579840 584942 580080 6 gpio_analog[5]
port 13 nsew signal bidirectional
rlabel metal3 s 583502 639272 584942 639512 6 gpio_analog[6]
port 14 nsew signal bidirectional
rlabel metal3 s -978 689592 462 689832 4 gpio_analog[7]
port 15 nsew signal bidirectional
rlabel metal3 s -978 670824 462 671064 4 gpio_analog[8]
port 16 nsew signal bidirectional
rlabel metal3 s -978 614520 462 614760 4 gpio_analog[9]
port 17 nsew signal bidirectional
rlabel metal3 s 583502 292336 584942 292576 6 gpio_noesd[0]
port 18 nsew signal bidirectional
rlabel metal3 s -978 548832 462 549072 4 gpio_noesd[10]
port 19 nsew signal bidirectional
rlabel metal3 s -978 492528 462 492768 4 gpio_noesd[11]
port 20 nsew signal bidirectional
rlabel metal3 s -978 436224 462 436464 4 gpio_noesd[12]
port 21 nsew signal bidirectional
rlabel metal3 s -978 379920 462 380160 4 gpio_noesd[13]
port 22 nsew signal bidirectional
rlabel metal3 s -978 323616 462 323856 4 gpio_noesd[14]
port 23 nsew signal bidirectional
rlabel metal3 s -978 267312 462 267552 4 gpio_noesd[15]
port 24 nsew signal bidirectional
rlabel metal3 s -978 211008 462 211248 4 gpio_noesd[16]
port 25 nsew signal bidirectional
rlabel metal3 s -978 154704 462 154944 4 gpio_noesd[17]
port 26 nsew signal bidirectional
rlabel metal3 s 583502 351768 584942 352008 6 gpio_noesd[1]
port 27 nsew signal bidirectional
rlabel metal3 s 583502 411200 584942 411440 6 gpio_noesd[2]
port 28 nsew signal bidirectional
rlabel metal3 s 583502 470768 584942 471008 6 gpio_noesd[3]
port 29 nsew signal bidirectional
rlabel metal3 s 583502 530200 584942 530440 6 gpio_noesd[4]
port 30 nsew signal bidirectional
rlabel metal3 s 583502 589768 584942 590008 6 gpio_noesd[5]
port 31 nsew signal bidirectional
rlabel metal3 s 583502 649200 584942 649440 6 gpio_noesd[6]
port 32 nsew signal bidirectional
rlabel metal3 s -978 680208 462 680448 4 gpio_noesd[7]
port 33 nsew signal bidirectional
rlabel metal3 s -978 661440 462 661680 4 gpio_noesd[8]
port 34 nsew signal bidirectional
rlabel metal3 s -978 605136 462 605376 4 gpio_noesd[9]
port 35 nsew signal bidirectional
rlabel metal3 s 583502 698840 584942 699080 6 io_analog[0]
port 36 nsew signal bidirectional
rlabel metal3 s -978 698976 462 699216 4 io_analog[10]
port 37 nsew signal bidirectional
rlabel metal2 s 564392 703508 564504 704948 6 io_analog[1]
port 38 nsew signal bidirectional
rlabel metal2 s 525476 703508 525588 704948 6 io_analog[2]
port 39 nsew signal bidirectional
rlabel metal2 s 486560 703508 486672 704948 6 io_analog[3]
port 40 nsew signal bidirectional
rlabel metal2 s 369720 703508 369832 704948 6 io_analog[4]
port 41 nsew signal bidirectional
rlabel metal2 s 252972 703508 253084 704948 6 io_analog[5]
port 42 nsew signal bidirectional
rlabel metal2 s 136132 703508 136244 704948 6 io_analog[6]
port 43 nsew signal bidirectional
rlabel metal2 s 97216 703508 97328 704948 6 io_analog[7]
port 44 nsew signal bidirectional
rlabel metal2 s 58300 703508 58412 704948 6 io_analog[8]
port 45 nsew signal bidirectional
rlabel metal2 s 19384 703508 19496 704948 6 io_analog[9]
port 46 nsew signal bidirectional
rlabel metal2 s 447644 703508 447756 704948 6 io_clamp_high[0]
port 47 nsew signal bidirectional
rlabel metal2 s 330804 703508 330916 704948 6 io_clamp_high[1]
port 48 nsew signal bidirectional
rlabel metal2 s 214056 703508 214168 704948 6 io_clamp_high[2]
port 49 nsew signal bidirectional
rlabel metal2 s 408728 703508 408840 704948 6 io_clamp_low[0]
port 50 nsew signal bidirectional
rlabel metal2 s 291888 703508 292000 704948 6 io_clamp_low[1]
port 51 nsew signal bidirectional
rlabel metal2 s 175048 703508 175160 704948 6 io_clamp_low[2]
port 52 nsew signal bidirectional
rlabel metal3 s 583502 14624 584942 14864 6 io_in[0]
port 53 nsew signal input
rlabel metal3 s 583502 24552 584942 24792 6 io_out[0]
port 54 nsew signal tristate
rlabel metal3 s 583502 490624 584942 490864 6 io_in[10]
port 55 nsew signal input
rlabel metal3 s 583502 500552 584942 500792 6 io_out[10]
port 56 nsew signal tristate
rlabel metal3 s 583502 550056 584942 550296 6 io_in[11]
port 57 nsew signal input
rlabel metal3 s 583502 559984 584942 560224 6 io_out[11]
port 58 nsew signal tristate
rlabel metal3 s 583502 609488 584942 609728 6 io_in[12]
port 59 nsew signal input
rlabel metal3 s 583502 619416 584942 619656 6 io_out[12]
port 60 nsew signal tristate
rlabel metal3 s 583502 669056 584942 669296 6 io_in[13]
port 61 nsew signal input
rlabel metal3 s 583502 678984 584942 679224 6 io_out[13]
port 62 nsew signal tristate
rlabel metal3 s -978 642672 462 642912 4 io_in[14]
port 63 nsew signal input
rlabel metal3 s -978 633288 462 633528 4 io_out[14]
port 64 nsew signal tristate
rlabel metal3 s -978 586368 462 586608 4 io_in[15]
port 65 nsew signal input
rlabel metal3 s -978 576984 462 577224 4 io_out[15]
port 66 nsew signal tristate
rlabel metal3 s -978 530064 462 530304 4 io_in[16]
port 67 nsew signal input
rlabel metal3 s -978 520680 462 520920 4 io_out[16]
port 68 nsew signal tristate
rlabel metal3 s -978 473760 462 474000 4 io_in[17]
port 69 nsew signal input
rlabel metal3 s -978 464376 462 464616 4 io_out[17]
port 70 nsew signal tristate
rlabel metal3 s -978 417456 462 417696 4 io_in[18]
port 71 nsew signal input
rlabel metal3 s -978 408072 462 408312 4 io_out[18]
port 72 nsew signal tristate
rlabel metal3 s -978 361152 462 361392 4 io_in[19]
port 73 nsew signal input
rlabel metal3 s -978 351768 462 352008 4 io_out[19]
port 74 nsew signal tristate
rlabel metal3 s 583502 54336 584942 54576 6 io_in[1]
port 75 nsew signal input
rlabel metal3 s 583502 64264 584942 64504 6 io_out[1]
port 76 nsew signal tristate
rlabel metal3 s -978 304848 462 305088 4 io_in[20]
port 77 nsew signal input
rlabel metal3 s -978 295464 462 295704 4 io_out[20]
port 78 nsew signal tristate
rlabel metal3 s -978 248544 462 248784 4 io_in[21]
port 79 nsew signal input
rlabel metal3 s -978 239160 462 239400 4 io_out[21]
port 80 nsew signal tristate
rlabel metal3 s -978 192240 462 192480 4 io_in[22]
port 81 nsew signal input
rlabel metal3 s -978 182856 462 183096 4 io_out[22]
port 82 nsew signal tristate
rlabel metal3 s -978 135936 462 136176 4 io_in[23]
port 83 nsew signal input
rlabel metal3 s -978 126552 462 126792 4 io_out[23]
port 84 nsew signal tristate
rlabel metal3 s -978 98400 462 98640 4 io_in[24]
port 85 nsew signal input
rlabel metal3 s -978 89016 462 89256 4 io_out[24]
port 86 nsew signal tristate
rlabel metal3 s -978 60864 462 61104 4 io_in[25]
port 87 nsew signal input
rlabel metal3 s -978 51480 462 51720 4 io_out[25]
port 88 nsew signal tristate
rlabel metal3 s -978 23328 462 23568 4 io_in[26]
port 89 nsew signal input
rlabel metal3 s -978 13944 462 14184 4 io_out[26]
port 90 nsew signal tristate
rlabel metal3 s 583502 94048 584942 94288 6 io_in[2]
port 91 nsew signal input
rlabel metal3 s 583502 103976 584942 104216 6 io_out[2]
port 92 nsew signal tristate
rlabel metal3 s 583502 133624 584942 133864 6 io_in[3]
port 93 nsew signal input
rlabel metal3 s 583502 143552 584942 143792 6 io_out[3]
port 94 nsew signal tristate
rlabel metal3 s 583502 173336 584942 173576 6 io_in[4]
port 95 nsew signal input
rlabel metal3 s 583502 183264 584942 183504 6 io_out[4]
port 96 nsew signal tristate
rlabel metal3 s 583502 212912 584942 213152 6 io_in[5]
port 97 nsew signal input
rlabel metal3 s 583502 222840 584942 223080 6 io_out[5]
port 98 nsew signal tristate
rlabel metal3 s 583502 252624 584942 252864 6 io_in[6]
port 99 nsew signal input
rlabel metal3 s 583502 262552 584942 262792 6 io_out[6]
port 100 nsew signal tristate
rlabel metal3 s 583502 312056 584942 312296 6 io_in[7]
port 101 nsew signal input
rlabel metal3 s 583502 321984 584942 322224 6 io_out[7]
port 102 nsew signal tristate
rlabel metal3 s 583502 371624 584942 371864 6 io_in[8]
port 103 nsew signal input
rlabel metal3 s 583502 381552 584942 381792 6 io_out[8]
port 104 nsew signal tristate
rlabel metal3 s 583502 431056 584942 431296 6 io_in[9]
port 105 nsew signal input
rlabel metal3 s 583502 440984 584942 441224 6 io_out[9]
port 106 nsew signal tristate
rlabel metal3 s 583502 4832 584942 5072 6 io_in_3v3[0]
port 107 nsew signal input
rlabel metal3 s 583502 480696 584942 480936 6 io_in_3v3[10]
port 108 nsew signal input
rlabel metal3 s 583502 540128 584942 540368 6 io_in_3v3[11]
port 109 nsew signal input
rlabel metal3 s 583502 599696 584942 599936 6 io_in_3v3[12]
port 110 nsew signal input
rlabel metal3 s 583502 659128 584942 659368 6 io_in_3v3[13]
port 111 nsew signal input
rlabel metal3 s -978 652056 462 652296 4 io_in_3v3[14]
port 112 nsew signal input
rlabel metal3 s -978 595752 462 595992 4 io_in_3v3[15]
port 113 nsew signal input
rlabel metal3 s -978 539448 462 539688 4 io_in_3v3[16]
port 114 nsew signal input
rlabel metal3 s -978 483144 462 483384 4 io_in_3v3[17]
port 115 nsew signal input
rlabel metal3 s -978 426840 462 427080 4 io_in_3v3[18]
port 116 nsew signal input
rlabel metal3 s -978 370536 462 370776 4 io_in_3v3[19]
port 117 nsew signal input
rlabel metal3 s 583502 44408 584942 44648 6 io_in_3v3[1]
port 118 nsew signal input
rlabel metal3 s -978 314232 462 314472 4 io_in_3v3[20]
port 119 nsew signal input
rlabel metal3 s -978 257928 462 258168 4 io_in_3v3[21]
port 120 nsew signal input
rlabel metal3 s -978 201624 462 201864 4 io_in_3v3[22]
port 121 nsew signal input
rlabel metal3 s -978 145320 462 145560 4 io_in_3v3[23]
port 122 nsew signal input
rlabel metal3 s -978 107784 462 108024 4 io_in_3v3[24]
port 123 nsew signal input
rlabel metal3 s -978 70248 462 70488 4 io_in_3v3[25]
port 124 nsew signal input
rlabel metal3 s -978 32712 462 32952 4 io_in_3v3[26]
port 125 nsew signal input
rlabel metal3 s 583502 84120 584942 84360 6 io_in_3v3[2]
port 126 nsew signal input
rlabel metal3 s 583502 123696 584942 123936 6 io_in_3v3[3]
port 127 nsew signal input
rlabel metal3 s 583502 163408 584942 163648 6 io_in_3v3[4]
port 128 nsew signal input
rlabel metal3 s 583502 203120 584942 203360 6 io_in_3v3[5]
port 129 nsew signal input
rlabel metal3 s 583502 242696 584942 242936 6 io_in_3v3[6]
port 130 nsew signal input
rlabel metal3 s 583502 302264 584942 302504 6 io_in_3v3[7]
port 131 nsew signal input
rlabel metal3 s 583502 361696 584942 361936 6 io_in_3v3[8]
port 132 nsew signal input
rlabel metal3 s 583502 421128 584942 421368 6 io_in_3v3[9]
port 133 nsew signal input
rlabel metal3 s 583502 34480 584942 34720 6 io_oeb[0]
port 134 nsew signal tristate
rlabel metal3 s 583502 510344 584942 510584 6 io_oeb[10]
port 135 nsew signal tristate
rlabel metal3 s 583502 569912 584942 570152 6 io_oeb[11]
port 136 nsew signal tristate
rlabel metal3 s 583502 629344 584942 629584 6 io_oeb[12]
port 137 nsew signal tristate
rlabel metal3 s 583502 688912 584942 689152 6 io_oeb[13]
port 138 nsew signal tristate
rlabel metal3 s -978 623904 462 624144 4 io_oeb[14]
port 139 nsew signal tristate
rlabel metal3 s -978 567600 462 567840 4 io_oeb[15]
port 140 nsew signal tristate
rlabel metal3 s -978 511296 462 511536 4 io_oeb[16]
port 141 nsew signal tristate
rlabel metal3 s -978 454992 462 455232 4 io_oeb[17]
port 142 nsew signal tristate
rlabel metal3 s -978 398688 462 398928 4 io_oeb[18]
port 143 nsew signal tristate
rlabel metal3 s -978 342384 462 342624 4 io_oeb[19]
port 144 nsew signal tristate
rlabel metal3 s 583502 74192 584942 74432 6 io_oeb[1]
port 145 nsew signal tristate
rlabel metal3 s -978 286080 462 286320 4 io_oeb[20]
port 146 nsew signal tristate
rlabel metal3 s -978 229776 462 230016 4 io_oeb[21]
port 147 nsew signal tristate
rlabel metal3 s -978 173472 462 173712 4 io_oeb[22]
port 148 nsew signal tristate
rlabel metal3 s -978 117168 462 117408 4 io_oeb[23]
port 149 nsew signal tristate
rlabel metal3 s -978 79632 462 79872 4 io_oeb[24]
port 150 nsew signal tristate
rlabel metal3 s -978 42096 462 42336 4 io_oeb[25]
port 151 nsew signal tristate
rlabel metal3 s -978 4560 462 4800 4 io_oeb[26]
port 152 nsew signal tristate
rlabel metal3 s 583502 113768 584942 114008 6 io_oeb[2]
port 153 nsew signal tristate
rlabel metal3 s 583502 153480 584942 153720 6 io_oeb[3]
port 154 nsew signal tristate
rlabel metal3 s 583502 193192 584942 193432 6 io_oeb[4]
port 155 nsew signal tristate
rlabel metal3 s 583502 232768 584942 233008 6 io_oeb[5]
port 156 nsew signal tristate
rlabel metal3 s 583502 272480 584942 272720 6 io_oeb[6]
port 157 nsew signal tristate
rlabel metal3 s 583502 331912 584942 332152 6 io_oeb[7]
port 158 nsew signal tristate
rlabel metal3 s 583502 391480 584942 391720 6 io_oeb[8]
port 159 nsew signal tristate
rlabel metal3 s 583502 450912 584942 451152 6 io_oeb[9]
port 160 nsew signal tristate
rlabel metal2 s 125828 -972 125940 468 8 la_data_in[0]
port 161 nsew signal input
rlabel metal2 s 480488 -972 480600 468 8 la_data_in[100]
port 162 nsew signal input
rlabel metal2 s 483984 -972 484096 468 8 la_data_in[101]
port 163 nsew signal input
rlabel metal2 s 487572 -972 487684 468 8 la_data_in[102]
port 164 nsew signal input
rlabel metal2 s 491068 -972 491180 468 8 la_data_in[103]
port 165 nsew signal input
rlabel metal2 s 494656 -972 494768 468 8 la_data_in[104]
port 166 nsew signal input
rlabel metal2 s 498152 -972 498264 468 8 la_data_in[105]
port 167 nsew signal input
rlabel metal2 s 501740 -972 501852 468 8 la_data_in[106]
port 168 nsew signal input
rlabel metal2 s 505328 -972 505440 468 8 la_data_in[107]
port 169 nsew signal input
rlabel metal2 s 508824 -972 508936 468 8 la_data_in[108]
port 170 nsew signal input
rlabel metal2 s 512412 -972 512524 468 8 la_data_in[109]
port 171 nsew signal input
rlabel metal2 s 161248 -972 161360 468 8 la_data_in[10]
port 172 nsew signal input
rlabel metal2 s 515908 -972 516020 468 8 la_data_in[110]
port 173 nsew signal input
rlabel metal2 s 519496 -972 519608 468 8 la_data_in[111]
port 174 nsew signal input
rlabel metal2 s 522992 -972 523104 468 8 la_data_in[112]
port 175 nsew signal input
rlabel metal2 s 526580 -972 526692 468 8 la_data_in[113]
port 176 nsew signal input
rlabel metal2 s 530076 -972 530188 468 8 la_data_in[114]
port 177 nsew signal input
rlabel metal2 s 533664 -972 533776 468 8 la_data_in[115]
port 178 nsew signal input
rlabel metal2 s 537160 -972 537272 468 8 la_data_in[116]
port 179 nsew signal input
rlabel metal2 s 540748 -972 540860 468 8 la_data_in[117]
port 180 nsew signal input
rlabel metal2 s 544336 -972 544448 468 8 la_data_in[118]
port 181 nsew signal input
rlabel metal2 s 547832 -972 547944 468 8 la_data_in[119]
port 182 nsew signal input
rlabel metal2 s 164836 -972 164948 468 8 la_data_in[11]
port 183 nsew signal input
rlabel metal2 s 551420 -972 551532 468 8 la_data_in[120]
port 184 nsew signal input
rlabel metal2 s 554916 -972 555028 468 8 la_data_in[121]
port 185 nsew signal input
rlabel metal2 s 558504 -972 558616 468 8 la_data_in[122]
port 186 nsew signal input
rlabel metal2 s 562000 -972 562112 468 8 la_data_in[123]
port 187 nsew signal input
rlabel metal2 s 565588 -972 565700 468 8 la_data_in[124]
port 188 nsew signal input
rlabel metal2 s 569084 -972 569196 468 8 la_data_in[125]
port 189 nsew signal input
rlabel metal2 s 572672 -972 572784 468 8 la_data_in[126]
port 190 nsew signal input
rlabel metal2 s 576260 -972 576372 468 8 la_data_in[127]
port 191 nsew signal input
rlabel metal2 s 168332 -972 168444 468 8 la_data_in[12]
port 192 nsew signal input
rlabel metal2 s 171920 -972 172032 468 8 la_data_in[13]
port 193 nsew signal input
rlabel metal2 s 175416 -972 175528 468 8 la_data_in[14]
port 194 nsew signal input
rlabel metal2 s 179004 -972 179116 468 8 la_data_in[15]
port 195 nsew signal input
rlabel metal2 s 182500 -972 182612 468 8 la_data_in[16]
port 196 nsew signal input
rlabel metal2 s 186088 -972 186200 468 8 la_data_in[17]
port 197 nsew signal input
rlabel metal2 s 189676 -972 189788 468 8 la_data_in[18]
port 198 nsew signal input
rlabel metal2 s 193172 -972 193284 468 8 la_data_in[19]
port 199 nsew signal input
rlabel metal2 s 129324 -972 129436 468 8 la_data_in[1]
port 200 nsew signal input
rlabel metal2 s 196760 -972 196872 468 8 la_data_in[20]
port 201 nsew signal input
rlabel metal2 s 200256 -972 200368 468 8 la_data_in[21]
port 202 nsew signal input
rlabel metal2 s 203844 -972 203956 468 8 la_data_in[22]
port 203 nsew signal input
rlabel metal2 s 207340 -972 207452 468 8 la_data_in[23]
port 204 nsew signal input
rlabel metal2 s 210928 -972 211040 468 8 la_data_in[24]
port 205 nsew signal input
rlabel metal2 s 214424 -972 214536 468 8 la_data_in[25]
port 206 nsew signal input
rlabel metal2 s 218012 -972 218124 468 8 la_data_in[26]
port 207 nsew signal input
rlabel metal2 s 221508 -972 221620 468 8 la_data_in[27]
port 208 nsew signal input
rlabel metal2 s 225096 -972 225208 468 8 la_data_in[28]
port 209 nsew signal input
rlabel metal2 s 228684 -972 228796 468 8 la_data_in[29]
port 210 nsew signal input
rlabel metal2 s 132912 -972 133024 468 8 la_data_in[2]
port 211 nsew signal input
rlabel metal2 s 232180 -972 232292 468 8 la_data_in[30]
port 212 nsew signal input
rlabel metal2 s 235768 -972 235880 468 8 la_data_in[31]
port 213 nsew signal input
rlabel metal2 s 239264 -972 239376 468 8 la_data_in[32]
port 214 nsew signal input
rlabel metal2 s 242852 -972 242964 468 8 la_data_in[33]
port 215 nsew signal input
rlabel metal2 s 246348 -972 246460 468 8 la_data_in[34]
port 216 nsew signal input
rlabel metal2 s 249936 -972 250048 468 8 la_data_in[35]
port 217 nsew signal input
rlabel metal2 s 253432 -972 253544 468 8 la_data_in[36]
port 218 nsew signal input
rlabel metal2 s 257020 -972 257132 468 8 la_data_in[37]
port 219 nsew signal input
rlabel metal2 s 260608 -972 260720 468 8 la_data_in[38]
port 220 nsew signal input
rlabel metal2 s 264104 -972 264216 468 8 la_data_in[39]
port 221 nsew signal input
rlabel metal2 s 136408 -972 136520 468 8 la_data_in[3]
port 222 nsew signal input
rlabel metal2 s 267692 -972 267804 468 8 la_data_in[40]
port 223 nsew signal input
rlabel metal2 s 271188 -972 271300 468 8 la_data_in[41]
port 224 nsew signal input
rlabel metal2 s 274776 -972 274888 468 8 la_data_in[42]
port 225 nsew signal input
rlabel metal2 s 278272 -972 278384 468 8 la_data_in[43]
port 226 nsew signal input
rlabel metal2 s 281860 -972 281972 468 8 la_data_in[44]
port 227 nsew signal input
rlabel metal2 s 285356 -972 285468 468 8 la_data_in[45]
port 228 nsew signal input
rlabel metal2 s 288944 -972 289056 468 8 la_data_in[46]
port 229 nsew signal input
rlabel metal2 s 292532 -972 292644 468 8 la_data_in[47]
port 230 nsew signal input
rlabel metal2 s 296028 -972 296140 468 8 la_data_in[48]
port 231 nsew signal input
rlabel metal2 s 299616 -972 299728 468 8 la_data_in[49]
port 232 nsew signal input
rlabel metal2 s 139996 -972 140108 468 8 la_data_in[4]
port 233 nsew signal input
rlabel metal2 s 303112 -972 303224 468 8 la_data_in[50]
port 234 nsew signal input
rlabel metal2 s 306700 -972 306812 468 8 la_data_in[51]
port 235 nsew signal input
rlabel metal2 s 310196 -972 310308 468 8 la_data_in[52]
port 236 nsew signal input
rlabel metal2 s 313784 -972 313896 468 8 la_data_in[53]
port 237 nsew signal input
rlabel metal2 s 317280 -972 317392 468 8 la_data_in[54]
port 238 nsew signal input
rlabel metal2 s 320868 -972 320980 468 8 la_data_in[55]
port 239 nsew signal input
rlabel metal2 s 324364 -972 324476 468 8 la_data_in[56]
port 240 nsew signal input
rlabel metal2 s 327952 -972 328064 468 8 la_data_in[57]
port 241 nsew signal input
rlabel metal2 s 331540 -972 331652 468 8 la_data_in[58]
port 242 nsew signal input
rlabel metal2 s 335036 -972 335148 468 8 la_data_in[59]
port 243 nsew signal input
rlabel metal2 s 143492 -972 143604 468 8 la_data_in[5]
port 244 nsew signal input
rlabel metal2 s 338624 -972 338736 468 8 la_data_in[60]
port 245 nsew signal input
rlabel metal2 s 342120 -972 342232 468 8 la_data_in[61]
port 246 nsew signal input
rlabel metal2 s 345708 -972 345820 468 8 la_data_in[62]
port 247 nsew signal input
rlabel metal2 s 349204 -972 349316 468 8 la_data_in[63]
port 248 nsew signal input
rlabel metal2 s 352792 -972 352904 468 8 la_data_in[64]
port 249 nsew signal input
rlabel metal2 s 356288 -972 356400 468 8 la_data_in[65]
port 250 nsew signal input
rlabel metal2 s 359876 -972 359988 468 8 la_data_in[66]
port 251 nsew signal input
rlabel metal2 s 363464 -972 363576 468 8 la_data_in[67]
port 252 nsew signal input
rlabel metal2 s 366960 -972 367072 468 8 la_data_in[68]
port 253 nsew signal input
rlabel metal2 s 370548 -972 370660 468 8 la_data_in[69]
port 254 nsew signal input
rlabel metal2 s 147080 -972 147192 468 8 la_data_in[6]
port 255 nsew signal input
rlabel metal2 s 374044 -972 374156 468 8 la_data_in[70]
port 256 nsew signal input
rlabel metal2 s 377632 -972 377744 468 8 la_data_in[71]
port 257 nsew signal input
rlabel metal2 s 381128 -972 381240 468 8 la_data_in[72]
port 258 nsew signal input
rlabel metal2 s 384716 -972 384828 468 8 la_data_in[73]
port 259 nsew signal input
rlabel metal2 s 388212 -972 388324 468 8 la_data_in[74]
port 260 nsew signal input
rlabel metal2 s 391800 -972 391912 468 8 la_data_in[75]
port 261 nsew signal input
rlabel metal2 s 395296 -972 395408 468 8 la_data_in[76]
port 262 nsew signal input
rlabel metal2 s 398884 -972 398996 468 8 la_data_in[77]
port 263 nsew signal input
rlabel metal2 s 402472 -972 402584 468 8 la_data_in[78]
port 264 nsew signal input
rlabel metal2 s 405968 -972 406080 468 8 la_data_in[79]
port 265 nsew signal input
rlabel metal2 s 150576 -972 150688 468 8 la_data_in[7]
port 266 nsew signal input
rlabel metal2 s 409556 -972 409668 468 8 la_data_in[80]
port 267 nsew signal input
rlabel metal2 s 413052 -972 413164 468 8 la_data_in[81]
port 268 nsew signal input
rlabel metal2 s 416640 -972 416752 468 8 la_data_in[82]
port 269 nsew signal input
rlabel metal2 s 420136 -972 420248 468 8 la_data_in[83]
port 270 nsew signal input
rlabel metal2 s 423724 -972 423836 468 8 la_data_in[84]
port 271 nsew signal input
rlabel metal2 s 427220 -972 427332 468 8 la_data_in[85]
port 272 nsew signal input
rlabel metal2 s 430808 -972 430920 468 8 la_data_in[86]
port 273 nsew signal input
rlabel metal2 s 434396 -972 434508 468 8 la_data_in[87]
port 274 nsew signal input
rlabel metal2 s 437892 -972 438004 468 8 la_data_in[88]
port 275 nsew signal input
rlabel metal2 s 441480 -972 441592 468 8 la_data_in[89]
port 276 nsew signal input
rlabel metal2 s 154164 -972 154276 468 8 la_data_in[8]
port 277 nsew signal input
rlabel metal2 s 444976 -972 445088 468 8 la_data_in[90]
port 278 nsew signal input
rlabel metal2 s 448564 -972 448676 468 8 la_data_in[91]
port 279 nsew signal input
rlabel metal2 s 452060 -972 452172 468 8 la_data_in[92]
port 280 nsew signal input
rlabel metal2 s 455648 -972 455760 468 8 la_data_in[93]
port 281 nsew signal input
rlabel metal2 s 459144 -972 459256 468 8 la_data_in[94]
port 282 nsew signal input
rlabel metal2 s 462732 -972 462844 468 8 la_data_in[95]
port 283 nsew signal input
rlabel metal2 s 466228 -972 466340 468 8 la_data_in[96]
port 284 nsew signal input
rlabel metal2 s 469816 -972 469928 468 8 la_data_in[97]
port 285 nsew signal input
rlabel metal2 s 473404 -972 473516 468 8 la_data_in[98]
port 286 nsew signal input
rlabel metal2 s 476900 -972 477012 468 8 la_data_in[99]
port 287 nsew signal input
rlabel metal2 s 157752 -972 157864 468 8 la_data_in[9]
port 288 nsew signal input
rlabel metal2 s 126932 -972 127044 468 8 la_data_out[0]
port 289 nsew signal tristate
rlabel metal2 s 481684 -972 481796 468 8 la_data_out[100]
port 290 nsew signal tristate
rlabel metal2 s 485180 -972 485292 468 8 la_data_out[101]
port 291 nsew signal tristate
rlabel metal2 s 488768 -972 488880 468 8 la_data_out[102]
port 292 nsew signal tristate
rlabel metal2 s 492264 -972 492376 468 8 la_data_out[103]
port 293 nsew signal tristate
rlabel metal2 s 495852 -972 495964 468 8 la_data_out[104]
port 294 nsew signal tristate
rlabel metal2 s 499348 -972 499460 468 8 la_data_out[105]
port 295 nsew signal tristate
rlabel metal2 s 502936 -972 503048 468 8 la_data_out[106]
port 296 nsew signal tristate
rlabel metal2 s 506432 -972 506544 468 8 la_data_out[107]
port 297 nsew signal tristate
rlabel metal2 s 510020 -972 510132 468 8 la_data_out[108]
port 298 nsew signal tristate
rlabel metal2 s 513516 -972 513628 468 8 la_data_out[109]
port 299 nsew signal tristate
rlabel metal2 s 162444 -972 162556 468 8 la_data_out[10]
port 300 nsew signal tristate
rlabel metal2 s 517104 -972 517216 468 8 la_data_out[110]
port 301 nsew signal tristate
rlabel metal2 s 520692 -972 520804 468 8 la_data_out[111]
port 302 nsew signal tristate
rlabel metal2 s 524188 -972 524300 468 8 la_data_out[112]
port 303 nsew signal tristate
rlabel metal2 s 527776 -972 527888 468 8 la_data_out[113]
port 304 nsew signal tristate
rlabel metal2 s 531272 -972 531384 468 8 la_data_out[114]
port 305 nsew signal tristate
rlabel metal2 s 534860 -972 534972 468 8 la_data_out[115]
port 306 nsew signal tristate
rlabel metal2 s 538356 -972 538468 468 8 la_data_out[116]
port 307 nsew signal tristate
rlabel metal2 s 541944 -972 542056 468 8 la_data_out[117]
port 308 nsew signal tristate
rlabel metal2 s 545440 -972 545552 468 8 la_data_out[118]
port 309 nsew signal tristate
rlabel metal2 s 549028 -972 549140 468 8 la_data_out[119]
port 310 nsew signal tristate
rlabel metal2 s 166032 -972 166144 468 8 la_data_out[11]
port 311 nsew signal tristate
rlabel metal2 s 552616 -972 552728 468 8 la_data_out[120]
port 312 nsew signal tristate
rlabel metal2 s 556112 -972 556224 468 8 la_data_out[121]
port 313 nsew signal tristate
rlabel metal2 s 559700 -972 559812 468 8 la_data_out[122]
port 314 nsew signal tristate
rlabel metal2 s 563196 -972 563308 468 8 la_data_out[123]
port 315 nsew signal tristate
rlabel metal2 s 566784 -972 566896 468 8 la_data_out[124]
port 316 nsew signal tristate
rlabel metal2 s 570280 -972 570392 468 8 la_data_out[125]
port 317 nsew signal tristate
rlabel metal2 s 573868 -972 573980 468 8 la_data_out[126]
port 318 nsew signal tristate
rlabel metal2 s 577364 -972 577476 468 8 la_data_out[127]
port 319 nsew signal tristate
rlabel metal2 s 169528 -972 169640 468 8 la_data_out[12]
port 320 nsew signal tristate
rlabel metal2 s 173116 -972 173228 468 8 la_data_out[13]
port 321 nsew signal tristate
rlabel metal2 s 176612 -972 176724 468 8 la_data_out[14]
port 322 nsew signal tristate
rlabel metal2 s 180200 -972 180312 468 8 la_data_out[15]
port 323 nsew signal tristate
rlabel metal2 s 183696 -972 183808 468 8 la_data_out[16]
port 324 nsew signal tristate
rlabel metal2 s 187284 -972 187396 468 8 la_data_out[17]
port 325 nsew signal tristate
rlabel metal2 s 190780 -972 190892 468 8 la_data_out[18]
port 326 nsew signal tristate
rlabel metal2 s 194368 -972 194480 468 8 la_data_out[19]
port 327 nsew signal tristate
rlabel metal2 s 130520 -972 130632 468 8 la_data_out[1]
port 328 nsew signal tristate
rlabel metal2 s 197864 -972 197976 468 8 la_data_out[20]
port 329 nsew signal tristate
rlabel metal2 s 201452 -972 201564 468 8 la_data_out[21]
port 330 nsew signal tristate
rlabel metal2 s 205040 -972 205152 468 8 la_data_out[22]
port 331 nsew signal tristate
rlabel metal2 s 208536 -972 208648 468 8 la_data_out[23]
port 332 nsew signal tristate
rlabel metal2 s 212124 -972 212236 468 8 la_data_out[24]
port 333 nsew signal tristate
rlabel metal2 s 215620 -972 215732 468 8 la_data_out[25]
port 334 nsew signal tristate
rlabel metal2 s 219208 -972 219320 468 8 la_data_out[26]
port 335 nsew signal tristate
rlabel metal2 s 222704 -972 222816 468 8 la_data_out[27]
port 336 nsew signal tristate
rlabel metal2 s 226292 -972 226404 468 8 la_data_out[28]
port 337 nsew signal tristate
rlabel metal2 s 229788 -972 229900 468 8 la_data_out[29]
port 338 nsew signal tristate
rlabel metal2 s 134108 -972 134220 468 8 la_data_out[2]
port 339 nsew signal tristate
rlabel metal2 s 233376 -972 233488 468 8 la_data_out[30]
port 340 nsew signal tristate
rlabel metal2 s 236964 -972 237076 468 8 la_data_out[31]
port 341 nsew signal tristate
rlabel metal2 s 240460 -972 240572 468 8 la_data_out[32]
port 342 nsew signal tristate
rlabel metal2 s 244048 -972 244160 468 8 la_data_out[33]
port 343 nsew signal tristate
rlabel metal2 s 247544 -972 247656 468 8 la_data_out[34]
port 344 nsew signal tristate
rlabel metal2 s 251132 -972 251244 468 8 la_data_out[35]
port 345 nsew signal tristate
rlabel metal2 s 254628 -972 254740 468 8 la_data_out[36]
port 346 nsew signal tristate
rlabel metal2 s 258216 -972 258328 468 8 la_data_out[37]
port 347 nsew signal tristate
rlabel metal2 s 261712 -972 261824 468 8 la_data_out[38]
port 348 nsew signal tristate
rlabel metal2 s 265300 -972 265412 468 8 la_data_out[39]
port 349 nsew signal tristate
rlabel metal2 s 137604 -972 137716 468 8 la_data_out[3]
port 350 nsew signal tristate
rlabel metal2 s 268796 -972 268908 468 8 la_data_out[40]
port 351 nsew signal tristate
rlabel metal2 s 272384 -972 272496 468 8 la_data_out[41]
port 352 nsew signal tristate
rlabel metal2 s 275972 -972 276084 468 8 la_data_out[42]
port 353 nsew signal tristate
rlabel metal2 s 279468 -972 279580 468 8 la_data_out[43]
port 354 nsew signal tristate
rlabel metal2 s 283056 -972 283168 468 8 la_data_out[44]
port 355 nsew signal tristate
rlabel metal2 s 286552 -972 286664 468 8 la_data_out[45]
port 356 nsew signal tristate
rlabel metal2 s 290140 -972 290252 468 8 la_data_out[46]
port 357 nsew signal tristate
rlabel metal2 s 293636 -972 293748 468 8 la_data_out[47]
port 358 nsew signal tristate
rlabel metal2 s 297224 -972 297336 468 8 la_data_out[48]
port 359 nsew signal tristate
rlabel metal2 s 300720 -972 300832 468 8 la_data_out[49]
port 360 nsew signal tristate
rlabel metal2 s 141192 -972 141304 468 8 la_data_out[4]
port 361 nsew signal tristate
rlabel metal2 s 304308 -972 304420 468 8 la_data_out[50]
port 362 nsew signal tristate
rlabel metal2 s 307896 -972 308008 468 8 la_data_out[51]
port 363 nsew signal tristate
rlabel metal2 s 311392 -972 311504 468 8 la_data_out[52]
port 364 nsew signal tristate
rlabel metal2 s 314980 -972 315092 468 8 la_data_out[53]
port 365 nsew signal tristate
rlabel metal2 s 318476 -972 318588 468 8 la_data_out[54]
port 366 nsew signal tristate
rlabel metal2 s 322064 -972 322176 468 8 la_data_out[55]
port 367 nsew signal tristate
rlabel metal2 s 325560 -972 325672 468 8 la_data_out[56]
port 368 nsew signal tristate
rlabel metal2 s 329148 -972 329260 468 8 la_data_out[57]
port 369 nsew signal tristate
rlabel metal2 s 332644 -972 332756 468 8 la_data_out[58]
port 370 nsew signal tristate
rlabel metal2 s 336232 -972 336344 468 8 la_data_out[59]
port 371 nsew signal tristate
rlabel metal2 s 144688 -972 144800 468 8 la_data_out[5]
port 372 nsew signal tristate
rlabel metal2 s 339820 -972 339932 468 8 la_data_out[60]
port 373 nsew signal tristate
rlabel metal2 s 343316 -972 343428 468 8 la_data_out[61]
port 374 nsew signal tristate
rlabel metal2 s 346904 -972 347016 468 8 la_data_out[62]
port 375 nsew signal tristate
rlabel metal2 s 350400 -972 350512 468 8 la_data_out[63]
port 376 nsew signal tristate
rlabel metal2 s 353988 -972 354100 468 8 la_data_out[64]
port 377 nsew signal tristate
rlabel metal2 s 357484 -972 357596 468 8 la_data_out[65]
port 378 nsew signal tristate
rlabel metal2 s 361072 -972 361184 468 8 la_data_out[66]
port 379 nsew signal tristate
rlabel metal2 s 364568 -972 364680 468 8 la_data_out[67]
port 380 nsew signal tristate
rlabel metal2 s 368156 -972 368268 468 8 la_data_out[68]
port 381 nsew signal tristate
rlabel metal2 s 371652 -972 371764 468 8 la_data_out[69]
port 382 nsew signal tristate
rlabel metal2 s 148276 -972 148388 468 8 la_data_out[6]
port 383 nsew signal tristate
rlabel metal2 s 375240 -972 375352 468 8 la_data_out[70]
port 384 nsew signal tristate
rlabel metal2 s 378828 -972 378940 468 8 la_data_out[71]
port 385 nsew signal tristate
rlabel metal2 s 382324 -972 382436 468 8 la_data_out[72]
port 386 nsew signal tristate
rlabel metal2 s 385912 -972 386024 468 8 la_data_out[73]
port 387 nsew signal tristate
rlabel metal2 s 389408 -972 389520 468 8 la_data_out[74]
port 388 nsew signal tristate
rlabel metal2 s 392996 -972 393108 468 8 la_data_out[75]
port 389 nsew signal tristate
rlabel metal2 s 396492 -972 396604 468 8 la_data_out[76]
port 390 nsew signal tristate
rlabel metal2 s 400080 -972 400192 468 8 la_data_out[77]
port 391 nsew signal tristate
rlabel metal2 s 403576 -972 403688 468 8 la_data_out[78]
port 392 nsew signal tristate
rlabel metal2 s 407164 -972 407276 468 8 la_data_out[79]
port 393 nsew signal tristate
rlabel metal2 s 151772 -972 151884 468 8 la_data_out[7]
port 394 nsew signal tristate
rlabel metal2 s 410752 -972 410864 468 8 la_data_out[80]
port 395 nsew signal tristate
rlabel metal2 s 414248 -972 414360 468 8 la_data_out[81]
port 396 nsew signal tristate
rlabel metal2 s 417836 -972 417948 468 8 la_data_out[82]
port 397 nsew signal tristate
rlabel metal2 s 421332 -972 421444 468 8 la_data_out[83]
port 398 nsew signal tristate
rlabel metal2 s 424920 -972 425032 468 8 la_data_out[84]
port 399 nsew signal tristate
rlabel metal2 s 428416 -972 428528 468 8 la_data_out[85]
port 400 nsew signal tristate
rlabel metal2 s 432004 -972 432116 468 8 la_data_out[86]
port 401 nsew signal tristate
rlabel metal2 s 435500 -972 435612 468 8 la_data_out[87]
port 402 nsew signal tristate
rlabel metal2 s 439088 -972 439200 468 8 la_data_out[88]
port 403 nsew signal tristate
rlabel metal2 s 442584 -972 442696 468 8 la_data_out[89]
port 404 nsew signal tristate
rlabel metal2 s 155360 -972 155472 468 8 la_data_out[8]
port 405 nsew signal tristate
rlabel metal2 s 446172 -972 446284 468 8 la_data_out[90]
port 406 nsew signal tristate
rlabel metal2 s 449760 -972 449872 468 8 la_data_out[91]
port 407 nsew signal tristate
rlabel metal2 s 453256 -972 453368 468 8 la_data_out[92]
port 408 nsew signal tristate
rlabel metal2 s 456844 -972 456956 468 8 la_data_out[93]
port 409 nsew signal tristate
rlabel metal2 s 460340 -972 460452 468 8 la_data_out[94]
port 410 nsew signal tristate
rlabel metal2 s 463928 -972 464040 468 8 la_data_out[95]
port 411 nsew signal tristate
rlabel metal2 s 467424 -972 467536 468 8 la_data_out[96]
port 412 nsew signal tristate
rlabel metal2 s 471012 -972 471124 468 8 la_data_out[97]
port 413 nsew signal tristate
rlabel metal2 s 474508 -972 474620 468 8 la_data_out[98]
port 414 nsew signal tristate
rlabel metal2 s 478096 -972 478208 468 8 la_data_out[99]
port 415 nsew signal tristate
rlabel metal2 s 158856 -972 158968 468 8 la_data_out[9]
port 416 nsew signal tristate
rlabel metal2 s 128128 -972 128240 468 8 la_oenb[0]
port 417 nsew signal input
rlabel metal2 s 482788 -972 482900 468 8 la_oenb[100]
port 418 nsew signal input
rlabel metal2 s 486376 -972 486488 468 8 la_oenb[101]
port 419 nsew signal input
rlabel metal2 s 489872 -972 489984 468 8 la_oenb[102]
port 420 nsew signal input
rlabel metal2 s 493460 -972 493572 468 8 la_oenb[103]
port 421 nsew signal input
rlabel metal2 s 497048 -972 497160 468 8 la_oenb[104]
port 422 nsew signal input
rlabel metal2 s 500544 -972 500656 468 8 la_oenb[105]
port 423 nsew signal input
rlabel metal2 s 504132 -972 504244 468 8 la_oenb[106]
port 424 nsew signal input
rlabel metal2 s 507628 -972 507740 468 8 la_oenb[107]
port 425 nsew signal input
rlabel metal2 s 511216 -972 511328 468 8 la_oenb[108]
port 426 nsew signal input
rlabel metal2 s 514712 -972 514824 468 8 la_oenb[109]
port 427 nsew signal input
rlabel metal2 s 163640 -972 163752 468 8 la_oenb[10]
port 428 nsew signal input
rlabel metal2 s 518300 -972 518412 468 8 la_oenb[110]
port 429 nsew signal input
rlabel metal2 s 521796 -972 521908 468 8 la_oenb[111]
port 430 nsew signal input
rlabel metal2 s 525384 -972 525496 468 8 la_oenb[112]
port 431 nsew signal input
rlabel metal2 s 528972 -972 529084 468 8 la_oenb[113]
port 432 nsew signal input
rlabel metal2 s 532468 -972 532580 468 8 la_oenb[114]
port 433 nsew signal input
rlabel metal2 s 536056 -972 536168 468 8 la_oenb[115]
port 434 nsew signal input
rlabel metal2 s 539552 -972 539664 468 8 la_oenb[116]
port 435 nsew signal input
rlabel metal2 s 543140 -972 543252 468 8 la_oenb[117]
port 436 nsew signal input
rlabel metal2 s 546636 -972 546748 468 8 la_oenb[118]
port 437 nsew signal input
rlabel metal2 s 550224 -972 550336 468 8 la_oenb[119]
port 438 nsew signal input
rlabel metal2 s 167136 -972 167248 468 8 la_oenb[11]
port 439 nsew signal input
rlabel metal2 s 553720 -972 553832 468 8 la_oenb[120]
port 440 nsew signal input
rlabel metal2 s 557308 -972 557420 468 8 la_oenb[121]
port 441 nsew signal input
rlabel metal2 s 560804 -972 560916 468 8 la_oenb[122]
port 442 nsew signal input
rlabel metal2 s 564392 -972 564504 468 8 la_oenb[123]
port 443 nsew signal input
rlabel metal2 s 567980 -972 568092 468 8 la_oenb[124]
port 444 nsew signal input
rlabel metal2 s 571476 -972 571588 468 8 la_oenb[125]
port 445 nsew signal input
rlabel metal2 s 575064 -972 575176 468 8 la_oenb[126]
port 446 nsew signal input
rlabel metal2 s 578560 -972 578672 468 8 la_oenb[127]
port 447 nsew signal input
rlabel metal2 s 170724 -972 170836 468 8 la_oenb[12]
port 448 nsew signal input
rlabel metal2 s 174220 -972 174332 468 8 la_oenb[13]
port 449 nsew signal input
rlabel metal2 s 177808 -972 177920 468 8 la_oenb[14]
port 450 nsew signal input
rlabel metal2 s 181396 -972 181508 468 8 la_oenb[15]
port 451 nsew signal input
rlabel metal2 s 184892 -972 185004 468 8 la_oenb[16]
port 452 nsew signal input
rlabel metal2 s 188480 -972 188592 468 8 la_oenb[17]
port 453 nsew signal input
rlabel metal2 s 191976 -972 192088 468 8 la_oenb[18]
port 454 nsew signal input
rlabel metal2 s 195564 -972 195676 468 8 la_oenb[19]
port 455 nsew signal input
rlabel metal2 s 131716 -972 131828 468 8 la_oenb[1]
port 456 nsew signal input
rlabel metal2 s 199060 -972 199172 468 8 la_oenb[20]
port 457 nsew signal input
rlabel metal2 s 202648 -972 202760 468 8 la_oenb[21]
port 458 nsew signal input
rlabel metal2 s 206144 -972 206256 468 8 la_oenb[22]
port 459 nsew signal input
rlabel metal2 s 209732 -972 209844 468 8 la_oenb[23]
port 460 nsew signal input
rlabel metal2 s 213320 -972 213432 468 8 la_oenb[24]
port 461 nsew signal input
rlabel metal2 s 216816 -972 216928 468 8 la_oenb[25]
port 462 nsew signal input
rlabel metal2 s 220404 -972 220516 468 8 la_oenb[26]
port 463 nsew signal input
rlabel metal2 s 223900 -972 224012 468 8 la_oenb[27]
port 464 nsew signal input
rlabel metal2 s 227488 -972 227600 468 8 la_oenb[28]
port 465 nsew signal input
rlabel metal2 s 230984 -972 231096 468 8 la_oenb[29]
port 466 nsew signal input
rlabel metal2 s 135212 -972 135324 468 8 la_oenb[2]
port 467 nsew signal input
rlabel metal2 s 234572 -972 234684 468 8 la_oenb[30]
port 468 nsew signal input
rlabel metal2 s 238068 -972 238180 468 8 la_oenb[31]
port 469 nsew signal input
rlabel metal2 s 241656 -972 241768 468 8 la_oenb[32]
port 470 nsew signal input
rlabel metal2 s 245152 -972 245264 468 8 la_oenb[33]
port 471 nsew signal input
rlabel metal2 s 248740 -972 248852 468 8 la_oenb[34]
port 472 nsew signal input
rlabel metal2 s 252328 -972 252440 468 8 la_oenb[35]
port 473 nsew signal input
rlabel metal2 s 255824 -972 255936 468 8 la_oenb[36]
port 474 nsew signal input
rlabel metal2 s 259412 -972 259524 468 8 la_oenb[37]
port 475 nsew signal input
rlabel metal2 s 262908 -972 263020 468 8 la_oenb[38]
port 476 nsew signal input
rlabel metal2 s 266496 -972 266608 468 8 la_oenb[39]
port 477 nsew signal input
rlabel metal2 s 138800 -972 138912 468 8 la_oenb[3]
port 478 nsew signal input
rlabel metal2 s 269992 -972 270104 468 8 la_oenb[40]
port 479 nsew signal input
rlabel metal2 s 273580 -972 273692 468 8 la_oenb[41]
port 480 nsew signal input
rlabel metal2 s 277076 -972 277188 468 8 la_oenb[42]
port 481 nsew signal input
rlabel metal2 s 280664 -972 280776 468 8 la_oenb[43]
port 482 nsew signal input
rlabel metal2 s 284252 -972 284364 468 8 la_oenb[44]
port 483 nsew signal input
rlabel metal2 s 287748 -972 287860 468 8 la_oenb[45]
port 484 nsew signal input
rlabel metal2 s 291336 -972 291448 468 8 la_oenb[46]
port 485 nsew signal input
rlabel metal2 s 294832 -972 294944 468 8 la_oenb[47]
port 486 nsew signal input
rlabel metal2 s 298420 -972 298532 468 8 la_oenb[48]
port 487 nsew signal input
rlabel metal2 s 301916 -972 302028 468 8 la_oenb[49]
port 488 nsew signal input
rlabel metal2 s 142388 -972 142500 468 8 la_oenb[4]
port 489 nsew signal input
rlabel metal2 s 305504 -972 305616 468 8 la_oenb[50]
port 490 nsew signal input
rlabel metal2 s 309000 -972 309112 468 8 la_oenb[51]
port 491 nsew signal input
rlabel metal2 s 312588 -972 312700 468 8 la_oenb[52]
port 492 nsew signal input
rlabel metal2 s 316176 -972 316288 468 8 la_oenb[53]
port 493 nsew signal input
rlabel metal2 s 319672 -972 319784 468 8 la_oenb[54]
port 494 nsew signal input
rlabel metal2 s 323260 -972 323372 468 8 la_oenb[55]
port 495 nsew signal input
rlabel metal2 s 326756 -972 326868 468 8 la_oenb[56]
port 496 nsew signal input
rlabel metal2 s 330344 -972 330456 468 8 la_oenb[57]
port 497 nsew signal input
rlabel metal2 s 333840 -972 333952 468 8 la_oenb[58]
port 498 nsew signal input
rlabel metal2 s 337428 -972 337540 468 8 la_oenb[59]
port 499 nsew signal input
rlabel metal2 s 145884 -972 145996 468 8 la_oenb[5]
port 500 nsew signal input
rlabel metal2 s 340924 -972 341036 468 8 la_oenb[60]
port 501 nsew signal input
rlabel metal2 s 344512 -972 344624 468 8 la_oenb[61]
port 502 nsew signal input
rlabel metal2 s 348008 -972 348120 468 8 la_oenb[62]
port 503 nsew signal input
rlabel metal2 s 351596 -972 351708 468 8 la_oenb[63]
port 504 nsew signal input
rlabel metal2 s 355184 -972 355296 468 8 la_oenb[64]
port 505 nsew signal input
rlabel metal2 s 358680 -972 358792 468 8 la_oenb[65]
port 506 nsew signal input
rlabel metal2 s 362268 -972 362380 468 8 la_oenb[66]
port 507 nsew signal input
rlabel metal2 s 365764 -972 365876 468 8 la_oenb[67]
port 508 nsew signal input
rlabel metal2 s 369352 -972 369464 468 8 la_oenb[68]
port 509 nsew signal input
rlabel metal2 s 372848 -972 372960 468 8 la_oenb[69]
port 510 nsew signal input
rlabel metal2 s 149472 -972 149584 468 8 la_oenb[6]
port 511 nsew signal input
rlabel metal2 s 376436 -972 376548 468 8 la_oenb[70]
port 512 nsew signal input
rlabel metal2 s 379932 -972 380044 468 8 la_oenb[71]
port 513 nsew signal input
rlabel metal2 s 383520 -972 383632 468 8 la_oenb[72]
port 514 nsew signal input
rlabel metal2 s 387108 -972 387220 468 8 la_oenb[73]
port 515 nsew signal input
rlabel metal2 s 390604 -972 390716 468 8 la_oenb[74]
port 516 nsew signal input
rlabel metal2 s 394192 -972 394304 468 8 la_oenb[75]
port 517 nsew signal input
rlabel metal2 s 397688 -972 397800 468 8 la_oenb[76]
port 518 nsew signal input
rlabel metal2 s 401276 -972 401388 468 8 la_oenb[77]
port 519 nsew signal input
rlabel metal2 s 404772 -972 404884 468 8 la_oenb[78]
port 520 nsew signal input
rlabel metal2 s 408360 -972 408472 468 8 la_oenb[79]
port 521 nsew signal input
rlabel metal2 s 152968 -972 153080 468 8 la_oenb[7]
port 522 nsew signal input
rlabel metal2 s 411856 -972 411968 468 8 la_oenb[80]
port 523 nsew signal input
rlabel metal2 s 415444 -972 415556 468 8 la_oenb[81]
port 524 nsew signal input
rlabel metal2 s 418940 -972 419052 468 8 la_oenb[82]
port 525 nsew signal input
rlabel metal2 s 422528 -972 422640 468 8 la_oenb[83]
port 526 nsew signal input
rlabel metal2 s 426116 -972 426228 468 8 la_oenb[84]
port 527 nsew signal input
rlabel metal2 s 429612 -972 429724 468 8 la_oenb[85]
port 528 nsew signal input
rlabel metal2 s 433200 -972 433312 468 8 la_oenb[86]
port 529 nsew signal input
rlabel metal2 s 436696 -972 436808 468 8 la_oenb[87]
port 530 nsew signal input
rlabel metal2 s 440284 -972 440396 468 8 la_oenb[88]
port 531 nsew signal input
rlabel metal2 s 443780 -972 443892 468 8 la_oenb[89]
port 532 nsew signal input
rlabel metal2 s 156556 -972 156668 468 8 la_oenb[8]
port 533 nsew signal input
rlabel metal2 s 447368 -972 447480 468 8 la_oenb[90]
port 534 nsew signal input
rlabel metal2 s 450864 -972 450976 468 8 la_oenb[91]
port 535 nsew signal input
rlabel metal2 s 454452 -972 454564 468 8 la_oenb[92]
port 536 nsew signal input
rlabel metal2 s 458040 -972 458152 468 8 la_oenb[93]
port 537 nsew signal input
rlabel metal2 s 461536 -972 461648 468 8 la_oenb[94]
port 538 nsew signal input
rlabel metal2 s 465124 -972 465236 468 8 la_oenb[95]
port 539 nsew signal input
rlabel metal2 s 468620 -972 468732 468 8 la_oenb[96]
port 540 nsew signal input
rlabel metal2 s 472208 -972 472320 468 8 la_oenb[97]
port 541 nsew signal input
rlabel metal2 s 475704 -972 475816 468 8 la_oenb[98]
port 542 nsew signal input
rlabel metal2 s 479292 -972 479404 468 8 la_oenb[99]
port 543 nsew signal input
rlabel metal2 s 160052 -972 160164 468 8 la_oenb[9]
port 544 nsew signal input
rlabel metal2 s 579756 -972 579868 468 8 user_clock2
port 545 nsew signal input
rlabel metal2 s 580952 -972 581064 468 8 user_irq[0]
port 546 nsew signal tristate
rlabel metal2 s 582148 -972 582260 468 8 user_irq[1]
port 547 nsew signal tristate
rlabel metal2 s 583344 -972 583456 468 8 user_irq[2]
port 548 nsew signal tristate
rlabel metal2 s 524 -972 636 468 8 wb_clk_i
port 549 nsew signal input
rlabel metal2 s 1628 -972 1740 468 8 wb_rst_i
port 550 nsew signal input
rlabel metal2 s 2824 -972 2936 468 8 wbs_ack_o
port 551 nsew signal tristate
rlabel metal2 s 7608 -972 7720 468 8 wbs_adr_i[0]
port 552 nsew signal input
rlabel metal2 s 47812 -972 47924 468 8 wbs_adr_i[10]
port 553 nsew signal input
rlabel metal2 s 51308 -972 51420 468 8 wbs_adr_i[11]
port 554 nsew signal input
rlabel metal2 s 54896 -972 55008 468 8 wbs_adr_i[12]
port 555 nsew signal input
rlabel metal2 s 58392 -972 58504 468 8 wbs_adr_i[13]
port 556 nsew signal input
rlabel metal2 s 61980 -972 62092 468 8 wbs_adr_i[14]
port 557 nsew signal input
rlabel metal2 s 65476 -972 65588 468 8 wbs_adr_i[15]
port 558 nsew signal input
rlabel metal2 s 69064 -972 69176 468 8 wbs_adr_i[16]
port 559 nsew signal input
rlabel metal2 s 72560 -972 72672 468 8 wbs_adr_i[17]
port 560 nsew signal input
rlabel metal2 s 76148 -972 76260 468 8 wbs_adr_i[18]
port 561 nsew signal input
rlabel metal2 s 79644 -972 79756 468 8 wbs_adr_i[19]
port 562 nsew signal input
rlabel metal2 s 12300 -972 12412 468 8 wbs_adr_i[1]
port 563 nsew signal input
rlabel metal2 s 83232 -972 83344 468 8 wbs_adr_i[20]
port 564 nsew signal input
rlabel metal2 s 86820 -972 86932 468 8 wbs_adr_i[21]
port 565 nsew signal input
rlabel metal2 s 90316 -972 90428 468 8 wbs_adr_i[22]
port 566 nsew signal input
rlabel metal2 s 93904 -972 94016 468 8 wbs_adr_i[23]
port 567 nsew signal input
rlabel metal2 s 97400 -972 97512 468 8 wbs_adr_i[24]
port 568 nsew signal input
rlabel metal2 s 100988 -972 101100 468 8 wbs_adr_i[25]
port 569 nsew signal input
rlabel metal2 s 104484 -972 104596 468 8 wbs_adr_i[26]
port 570 nsew signal input
rlabel metal2 s 108072 -972 108184 468 8 wbs_adr_i[27]
port 571 nsew signal input
rlabel metal2 s 111568 -972 111680 468 8 wbs_adr_i[28]
port 572 nsew signal input
rlabel metal2 s 115156 -972 115268 468 8 wbs_adr_i[29]
port 573 nsew signal input
rlabel metal2 s 16992 -972 17104 468 8 wbs_adr_i[2]
port 574 nsew signal input
rlabel metal2 s 118744 -972 118856 468 8 wbs_adr_i[30]
port 575 nsew signal input
rlabel metal2 s 122240 -972 122352 468 8 wbs_adr_i[31]
port 576 nsew signal input
rlabel metal2 s 21776 -972 21888 468 8 wbs_adr_i[3]
port 577 nsew signal input
rlabel metal2 s 26468 -972 26580 468 8 wbs_adr_i[4]
port 578 nsew signal input
rlabel metal2 s 30056 -972 30168 468 8 wbs_adr_i[5]
port 579 nsew signal input
rlabel metal2 s 33552 -972 33664 468 8 wbs_adr_i[6]
port 580 nsew signal input
rlabel metal2 s 37140 -972 37252 468 8 wbs_adr_i[7]
port 581 nsew signal input
rlabel metal2 s 40636 -972 40748 468 8 wbs_adr_i[8]
port 582 nsew signal input
rlabel metal2 s 44224 -972 44336 468 8 wbs_adr_i[9]
port 583 nsew signal input
rlabel metal2 s 4020 -972 4132 468 8 wbs_cyc_i
port 584 nsew signal input
rlabel metal2 s 8712 -972 8824 468 8 wbs_dat_i[0]
port 585 nsew signal input
rlabel metal2 s 48916 -972 49028 468 8 wbs_dat_i[10]
port 586 nsew signal input
rlabel metal2 s 52504 -972 52616 468 8 wbs_dat_i[11]
port 587 nsew signal input
rlabel metal2 s 56000 -972 56112 468 8 wbs_dat_i[12]
port 588 nsew signal input
rlabel metal2 s 59588 -972 59700 468 8 wbs_dat_i[13]
port 589 nsew signal input
rlabel metal2 s 63176 -972 63288 468 8 wbs_dat_i[14]
port 590 nsew signal input
rlabel metal2 s 66672 -972 66784 468 8 wbs_dat_i[15]
port 591 nsew signal input
rlabel metal2 s 70260 -972 70372 468 8 wbs_dat_i[16]
port 592 nsew signal input
rlabel metal2 s 73756 -972 73868 468 8 wbs_dat_i[17]
port 593 nsew signal input
rlabel metal2 s 77344 -972 77456 468 8 wbs_dat_i[18]
port 594 nsew signal input
rlabel metal2 s 80840 -972 80952 468 8 wbs_dat_i[19]
port 595 nsew signal input
rlabel metal2 s 13496 -972 13608 468 8 wbs_dat_i[1]
port 596 nsew signal input
rlabel metal2 s 84428 -972 84540 468 8 wbs_dat_i[20]
port 597 nsew signal input
rlabel metal2 s 87924 -972 88036 468 8 wbs_dat_i[21]
port 598 nsew signal input
rlabel metal2 s 91512 -972 91624 468 8 wbs_dat_i[22]
port 599 nsew signal input
rlabel metal2 s 95100 -972 95212 468 8 wbs_dat_i[23]
port 600 nsew signal input
rlabel metal2 s 98596 -972 98708 468 8 wbs_dat_i[24]
port 601 nsew signal input
rlabel metal2 s 102184 -972 102296 468 8 wbs_dat_i[25]
port 602 nsew signal input
rlabel metal2 s 105680 -972 105792 468 8 wbs_dat_i[26]
port 603 nsew signal input
rlabel metal2 s 109268 -972 109380 468 8 wbs_dat_i[27]
port 604 nsew signal input
rlabel metal2 s 112764 -972 112876 468 8 wbs_dat_i[28]
port 605 nsew signal input
rlabel metal2 s 116352 -972 116464 468 8 wbs_dat_i[29]
port 606 nsew signal input
rlabel metal2 s 18188 -972 18300 468 8 wbs_dat_i[2]
port 607 nsew signal input
rlabel metal2 s 119848 -972 119960 468 8 wbs_dat_i[30]
port 608 nsew signal input
rlabel metal2 s 123436 -972 123548 468 8 wbs_dat_i[31]
port 609 nsew signal input
rlabel metal2 s 22972 -972 23084 468 8 wbs_dat_i[3]
port 610 nsew signal input
rlabel metal2 s 27664 -972 27776 468 8 wbs_dat_i[4]
port 611 nsew signal input
rlabel metal2 s 31252 -972 31364 468 8 wbs_dat_i[5]
port 612 nsew signal input
rlabel metal2 s 34748 -972 34860 468 8 wbs_dat_i[6]
port 613 nsew signal input
rlabel metal2 s 38336 -972 38448 468 8 wbs_dat_i[7]
port 614 nsew signal input
rlabel metal2 s 41832 -972 41944 468 8 wbs_dat_i[8]
port 615 nsew signal input
rlabel metal2 s 45420 -972 45532 468 8 wbs_dat_i[9]
port 616 nsew signal input
rlabel metal2 s 9908 -972 10020 468 8 wbs_dat_o[0]
port 617 nsew signal tristate
rlabel metal2 s 50112 -972 50224 468 8 wbs_dat_o[10]
port 618 nsew signal tristate
rlabel metal2 s 53700 -972 53812 468 8 wbs_dat_o[11]
port 619 nsew signal tristate
rlabel metal2 s 57196 -972 57308 468 8 wbs_dat_o[12]
port 620 nsew signal tristate
rlabel metal2 s 60784 -972 60896 468 8 wbs_dat_o[13]
port 621 nsew signal tristate
rlabel metal2 s 64280 -972 64392 468 8 wbs_dat_o[14]
port 622 nsew signal tristate
rlabel metal2 s 67868 -972 67980 468 8 wbs_dat_o[15]
port 623 nsew signal tristate
rlabel metal2 s 71456 -972 71568 468 8 wbs_dat_o[16]
port 624 nsew signal tristate
rlabel metal2 s 74952 -972 75064 468 8 wbs_dat_o[17]
port 625 nsew signal tristate
rlabel metal2 s 78540 -972 78652 468 8 wbs_dat_o[18]
port 626 nsew signal tristate
rlabel metal2 s 82036 -972 82148 468 8 wbs_dat_o[19]
port 627 nsew signal tristate
rlabel metal2 s 14692 -972 14804 468 8 wbs_dat_o[1]
port 628 nsew signal tristate
rlabel metal2 s 85624 -972 85736 468 8 wbs_dat_o[20]
port 629 nsew signal tristate
rlabel metal2 s 89120 -972 89232 468 8 wbs_dat_o[21]
port 630 nsew signal tristate
rlabel metal2 s 92708 -972 92820 468 8 wbs_dat_o[22]
port 631 nsew signal tristate
rlabel metal2 s 96204 -972 96316 468 8 wbs_dat_o[23]
port 632 nsew signal tristate
rlabel metal2 s 99792 -972 99904 468 8 wbs_dat_o[24]
port 633 nsew signal tristate
rlabel metal2 s 103288 -972 103400 468 8 wbs_dat_o[25]
port 634 nsew signal tristate
rlabel metal2 s 106876 -972 106988 468 8 wbs_dat_o[26]
port 635 nsew signal tristate
rlabel metal2 s 110464 -972 110576 468 8 wbs_dat_o[27]
port 636 nsew signal tristate
rlabel metal2 s 113960 -972 114072 468 8 wbs_dat_o[28]
port 637 nsew signal tristate
rlabel metal2 s 117548 -972 117660 468 8 wbs_dat_o[29]
port 638 nsew signal tristate
rlabel metal2 s 19384 -972 19496 468 8 wbs_dat_o[2]
port 639 nsew signal tristate
rlabel metal2 s 121044 -972 121156 468 8 wbs_dat_o[30]
port 640 nsew signal tristate
rlabel metal2 s 124632 -972 124744 468 8 wbs_dat_o[31]
port 641 nsew signal tristate
rlabel metal2 s 24168 -972 24280 468 8 wbs_dat_o[3]
port 642 nsew signal tristate
rlabel metal2 s 28860 -972 28972 468 8 wbs_dat_o[4]
port 643 nsew signal tristate
rlabel metal2 s 32356 -972 32468 468 8 wbs_dat_o[5]
port 644 nsew signal tristate
rlabel metal2 s 35944 -972 36056 468 8 wbs_dat_o[6]
port 645 nsew signal tristate
rlabel metal2 s 39532 -972 39644 468 8 wbs_dat_o[7]
port 646 nsew signal tristate
rlabel metal2 s 43028 -972 43140 468 8 wbs_dat_o[8]
port 647 nsew signal tristate
rlabel metal2 s 46616 -972 46728 468 8 wbs_dat_o[9]
port 648 nsew signal tristate
rlabel metal2 s 11104 -972 11216 468 8 wbs_sel_i[0]
port 649 nsew signal input
rlabel metal2 s 15888 -972 16000 468 8 wbs_sel_i[1]
port 650 nsew signal input
rlabel metal2 s 20580 -972 20692 468 8 wbs_sel_i[2]
port 651 nsew signal input
rlabel metal2 s 25272 -972 25384 468 8 wbs_sel_i[3]
port 652 nsew signal input
rlabel metal2 s 5216 -972 5328 468 8 wbs_stb_i
port 653 nsew signal input
rlabel metal2 s 6412 -972 6524 468 8 wbs_we_i
port 654 nsew signal input
rlabel metal4 s 585302 -936 585902 704848 6 vccd1
port 655 nsew power bidirectional
rlabel metal4 s -2014 -936 -1414 704848 4 vccd1.extra1
port 656 nsew power bidirectional
rlabel metal5 s -2014 704248 585902 704848 6 vccd1.extra2
port 657 nsew power bidirectional
rlabel metal5 s -2014 -936 585902 -336 8 vccd1.extra3
port 658 nsew power bidirectional
rlabel metal4 s 586242 -1876 586842 705788 6 vssd1
port 659 nsew ground bidirectional
rlabel metal4 s -2954 -1876 -2354 705788 4 vssd1.extra1
port 660 nsew ground bidirectional
rlabel metal5 s -2954 705188 586842 705788 6 vssd1.extra2
port 661 nsew ground bidirectional
rlabel metal5 s -2954 -1876 586842 -1276 8 vssd1.extra3
port 662 nsew ground bidirectional
rlabel metal4 s 587182 -2816 587782 706728 6 vccd2
port 663 nsew power bidirectional
rlabel metal4 s -3894 -2816 -3294 706728 4 vccd2.extra1
port 664 nsew power bidirectional
rlabel metal5 s -3894 706128 587782 706728 6 vccd2.extra2
port 665 nsew power bidirectional
rlabel metal5 s -3894 -2816 587782 -2216 8 vccd2.extra3
port 666 nsew power bidirectional
rlabel metal4 s 588122 -3756 588722 707668 6 vssd2
port 667 nsew ground bidirectional
rlabel metal4 s -4834 -3756 -4234 707668 4 vssd2.extra1
port 668 nsew ground bidirectional
rlabel metal5 s -4834 707068 588722 707668 6 vssd2.extra2
port 669 nsew ground bidirectional
rlabel metal5 s -4834 -3756 588722 -3156 8 vssd2.extra3
port 670 nsew ground bidirectional
rlabel metal4 s 589062 -4696 589662 708608 6 vdda1
port 671 nsew power bidirectional
rlabel metal4 s -5774 -4696 -5174 708608 4 vdda1.extra1
port 672 nsew power bidirectional
rlabel metal5 s -5774 708008 589662 708608 6 vdda1.extra2
port 673 nsew power bidirectional
rlabel metal5 s -5774 -4696 589662 -4096 8 vdda1.extra3
port 674 nsew power bidirectional
rlabel metal4 s 590002 -5636 590602 709548 6 vssa1
port 675 nsew ground bidirectional
rlabel metal4 s -6714 -5636 -6114 709548 4 vssa1.extra1
port 676 nsew ground bidirectional
rlabel metal5 s -6714 708948 590602 709548 6 vssa1.extra2
port 677 nsew ground bidirectional
rlabel metal5 s -6714 -5636 590602 -5036 8 vssa1.extra3
port 678 nsew ground bidirectional
rlabel metal4 s 590942 -6576 591542 710488 6 vdda2
port 679 nsew power bidirectional
rlabel metal4 s -7654 -6576 -7054 710488 4 vdda2.extra1
port 680 nsew power bidirectional
rlabel metal5 s -7654 709888 591542 710488 6 vdda2.extra2
port 681 nsew power bidirectional
rlabel metal5 s -7654 -6576 591542 -5976 8 vdda2.extra3
port 682 nsew power bidirectional
rlabel metal4 s 591882 -7516 592482 711428 6 vssa2
port 683 nsew ground bidirectional
rlabel metal4 s -8594 -7516 -7994 711428 4 vssa2.extra1
port 684 nsew ground bidirectional
rlabel metal5 s -8594 710828 592482 711428 6 vssa2.extra2
port 685 nsew ground bidirectional
rlabel metal5 s -8594 -7516 592482 -6916 8 vssa2.extra3
port 686 nsew ground bidirectional
<< end >>
