magic
tech sky130A
magscale 1 2
timestamp 1619633287
use user_analog_proj_example  user_analog_proj_example_0
timestamp 1619633287
transform 1 0 264772 0 1 616578
box -59 -22 25476 8324
use user_analog_project_wrapper_empty  user_analog_project_wrapper_empty_0
timestamp 1619448499
transform 1 0 -18 0 1 -12
box -8576 -7506 592500 711442
<< end >>
