  X �     0�     0 LIB  >A�7KƧ�9D�/��ZT �     0�     0 $$$CONTEXT_INFO$$$ 
  via_new           +  ,PCELL=via_new  +  ,P(width)=##0.25  +  ,P(starting_metal)=#l-4 +  ,P(length)=##0.5  +  ,P(hv)=false  +  ,P(ending_metal)=#l0  +   ,LIB=SKY130   
  mimcap_1          +  ,PCELL=mimcap_1 +  ,P(y_spacing)=##1 +  ,P(x_spacing)=##1 +  ,P(w)=##15  +  ,P(totalcap)=##450  +  ,P(l)=##15  +  ,P(array_y)=#l1 +  ,P(array_x)=#l1 +   ,LIB=SKY130   
  via_new$1           +  ,PCELL=via_new  +  ,P(width)=##0.48  +  ,P(starting_metal)=#l0  +  ,P(length)=##3  +  ,P(hv)=false  +  ,P(ending_metal)=#l3  +   ,LIB=SKY130   
  via_new$3           +  ,PCELL=via_new  +  ,P(width)=##5 +  ,P(starting_metal)=#l0  +  ,P(length)=##2  +  ,P(hv)=false  +  ,P(ending_metal)=#l3  +   ,LIB=SKY130   
  via_new$4           +  ,PCELL=via_new  +  ,P(width)=##0.4 +  ,P(starting_metal)=#l-1 +  ,P(length)=##2  +  ,P(hv)=false  +  ,P(ending_metal)=#l0  +   ,LIB=SKY130     �     0�     0 via_new  	   B   !     �           �       	   _   !     � ����      X       	   C   !      �           �       	   D   !      �           �          C  , ,   �����   �   U  O   U  O����   �����     �     0�     0 *sky130_fd_pr__res_xhigh_po_0p69_GF6QJT   �     0�     0 "sky130_fd_pr__pfet_01v8_VCXY4W    B   ,  6����<  6�    8;    8;���<  6����<      B   ,  6�  �  6�  
F  8;  
F  8;  �  6�  �      B   ,  6�    6�  f  8;  f  8;    6�        B   ,  6�  \  6�  �  8;  �  8;  \  6�  \      B   ,  6�����  6�   �  8;   �  8;����  6�����      B   ,  6�����  6����&  8;���&  8;����  6�����      B   ,  6����  6����f  8;���f  8;���  6����      B   ,  .    .  �  6�  �  6�    .        B   ,  .  6  .  �  6�  �  6�  6  .  6      B   ,  .  	V  .  	�  6�  	�  6�  	V  .  	V      B   ,  .  v  .    6�    6�  v  .  v      B   ,  .  �  .  ,  6�  ,  6�  �  .  �      B   ,  .  �  .  L  6�  L  6�  �  .  �      B   ,  .  �  .  l  6�  l  6�  �  .  �      B   ,  .����  .   �  6�   �  6�����  .����      B   ,  .���  .����  6�����  6����  .���      B   ,  .���6  .����  6�����  6����6  .���6      B   ,  .���V  .����  6�����  6����V  .���V      B   ,  .���v  .���  6����  6����v  .���v      B   ,  .����  .���,  6����,  6�����  .����      B   ,  6�  �  6�    8;    8;  �  6�  �      B   ,  6�  
�  6�  &  8;  &  8;  
�  6�  
�      B   ,  6�  <  6�  �  8;  �  8;  <  6�  <      B   ,  6�  |  6�  �  8;  �  8;  |  6�  |      B   ,  6�����  6����  8;���  8;����  6�����      B   ,  6�����  6����F  8;���F  8;����  6�����      B   ,  6����<  6�����  8;����  8;���<  6����<      _   ,  6����(  6�    8O    8O���(  6����(      C   ,  *����b  *�  �  +�  �  +����b  *����b      C   ,  +�  6  +�  �  9?  �  9?  6  +�  6      C   ,  7A  
�  7A  &  7�  &  7�  
�  7A  
�      C   ,  7A    7A  f  7�  f  7�    7A        C   ,  7A  \  7A  �  7�  �  7�  \  7A  \      C   ,  7A����  7A   �  7�   �  7�����  7A����      C   ,  7A����  7A���&  7����&  7�����  7A����      C   ,  7A���  7A���f  7����f  7����  7A���      C   ,  .r  �  .r  �  6j  �  6j  �  .r  �      C   ,  .r    .r  �  6j  �  6j    .r        C   ,  .r  
<  .r  
�  6j  
�  6j  
<  .r  
<      C   ,  .r  \  .r  	  6j  	  6j  \  .r  \      C   ,  .r  |  .r  &  6j  &  6j  |  .r  |      C   ,  .r  �  .r  F  6j  F  6j  �  .r  �      C   ,  .r  �  .r  f  6j  f  6j  �  .r  �      C   ,  .r   �  .r  �  6j  �  6j   �  .r   �      C   ,  .r����  .r����  6j����  6j����  .r����      C   ,  .r���  .r����  6j����  6j���  .r���      C   ,  .r���<  .r����  6j����  6j���<  .r���<      C   ,  .r���\  .r���  6j���  6j���\  .r���\      C   ,  .r���|  .r���&  6j���&  6j���|  .r���|      C   ,  .r����  .r���F  6j���F  6j����  .r����      C   ,  7A  �  7A    7�    7�  �  7A  �      C   ,  7A  �  7A  
F  7�  
F  7�  �  7A  �      C   ,  7A  <  7A  �  7�  �  7�  <  7A  <      C   ,  7A  |  7A  �  7�  �  7�  |  7A  |      C   ,  7A����  7A���  7����  7�����  7A����      C   ,  7A����  7A���F  7����F  7�����  7A����      C   ,  7A���<  7A����  7�����  7����<  7A���<      C   ,  +����b  +����  9?���  9?���b  +����b      C   ,  9?���b  9?  �  9�  �  9����b  9?���b      C   ,  7A���<  7A    7�    7����<  7A���<      D   ,  7#  
�  7#    8	    8	  
�  7#  
�      D   ,  7#  0  7#  R  8	  R  8	  0  7#  0      D   ,  7#  p  7#  �  8	  �  8	  p  7#  p      D   ,  7#����  7#   �  8	   �  8	����  7#����      D   ,  7#����  7#���  8	���  8	����  7#����      D   ,  7#���0  7#���R  8	���R  8	���0  7#���0      D   ,  .�  
  .�    6V    6V  
  .�  
      D   ,  ,[  >  ,[  	$  4+  	$  4+  >  ,[  >      D   ,  .�  ^  .�  D  6V  D  6V  ^  .�  ^      D   ,  ,[  ~  ,[  d  4+  d  4+  ~  ,[  ~      D   ,  .�  �  .�  �  6V  �  6V  �  .�  �      D   ,  ,[   �  ,[  �  4+  �  4+   �  ,[   �      D   ,  .�����  .�����  6V����  6V����  .�����      D   ,  ,[����  ,[����  4+����  4+����  ,[����      D   ,  .����  .����  6V���  6V���  .����      D   ,  ,[���>  ,[���$  4+���$  4+���>  ,[���>      D   ,  .����^  .����D  6V���D  6V���^  .����^      D   ,  .����~  .����d  6V���d  6V���~  .����~      D   ,  7#  �  7#  �  8	  �  8	  �  7#  �      D   ,  7#  	  7#  
2  8	  
2  8	  	  7#  	      D   ,  7#  P  7#  r  8	  r  8	  P  7#  P      D   ,  7#  �  7#  �  8	  �  8	  �  7#  �      D   ,  7#����  7#����  8	����  8	����  7#����      D   ,  7#���  7#���2  8	���2  8	���  7#���      D   ,  7#���P  7#���r  8	���r  8	���P  7#���P      D   ,  7#���P  7#  �  8�  �  8����P  7#���P      D   ,  ,[  �  ,[  �  4+  �  4+  �  ,[  �      D   ,  ,[  �  ,[  �  4+  �  4+  �  ,[  �      C  , ,  2���\  2���  2����  2����\  2���\      C  , ,  2���|  2���&  2����&  2����|  2���|      C  , ,  2����  2���F  2����F  2�����  2����      C  , ,  3�  
<  3�  
�  4+  
�  4+  
<  3�  
<      C  , ,  3�  |  3�  &  4+  &  4+  |  3�  |      C  , ,  3�  �  3�  f  4+  f  4+  �  3�  �      C  , ,  3�����  3�����  4+����  4+����  3�����      C  , ,  3����<  3�����  4+����  4+���<  3����<      C  , ,  3����|  3����&  4+���&  4+���|  3����|      C  , ,  3�����  3����F  4+���F  4+����  3�����      C  , ,  4�  
<  4�  
�  5�  
�  5�  
<  4�  
<      C  , ,  4�  |  4�  &  5�  &  5�  |  4�  |      C  , ,  4�  �  4�  f  5�  f  5�  �  4�  �      C  , ,  4�����  4�����  5�����  5�����  4�����      C  , ,  4����<  4�����  5�����  5����<  4����<      C  , ,  4����|  4����&  5����&  5����|  4����|      C  , ,  4�����  4����F  5����F  5�����  4�����      C  , ,  7A    7A  �  7�  �  7�    7A        C  , ,  7A  	L  7A  	�  7�  	�  7�  	L  7A  	L      C  , ,  7A  �  7A  6  7�  6  7�  �  7A  �      C  , ,  7A  �  7A  v  7�  v  7�  �  7A  �      C  , ,  7A���  7A����  7�����  7����  7A���      C  , ,  7A���L  7A����  7�����  7����L  7A���L      C  , ,  7A����  7A���6  7����6  7�����  7A����      C  , ,  7A  ,  7A  �  7�  �  7�  ,  7A  ,      C  , ,  7A  l  7A    7�    7�  l  7A  l      C  , ,  7A  �  7A  V  7�  V  7�  �  7A  �      C  , ,  7A����  7A   �  7�   �  7�����  7A����      C  , ,  7A���,  7A����  7�����  7����,  7A���,      C  , ,  7A���l  7A���  7����  7����l  7A���l      C  , ,  /I  �  /I  �  /�  �  /�  �  /I  �      C  , ,  /I    /I  �  /�  �  /�    /I        C  , ,  /I  
<  /I  
�  /�  
�  /�  
<  /I  
<      C  , ,  /I  \  /I  	  /�  	  /�  \  /I  \      C  , ,  /I  |  /I  &  /�  &  /�  |  /I  |      C  , ,  /I  �  /I  F  /�  F  /�  �  /I  �      C  , ,  /I  �  /I  f  /�  f  /�  �  /I  �      C  , ,  /I   �  /I  �  /�  �  /�   �  /I   �      C  , ,  /I����  /I����  /�����  /�����  /I����      C  , ,  /I���  /I����  /�����  /����  /I���      C  , ,  /I���<  /I����  /�����  /����<  /I���<      C  , ,  /I���\  /I���  /����  /����\  /I���\      C  , ,  /I���|  /I���&  /����&  /����|  /I���|      C  , ,  /I����  /I���F  /����F  /�����  /I����      C  , ,  0�  �  0�  �  1[  �  1[  �  0�  �      C  , ,  0�    0�  �  1[  �  1[    0�        C  , ,  0�  
<  0�  
�  1[  
�  1[  
<  0�  
<      C  , ,  0�  \  0�  	  1[  	  1[  \  0�  \      C  , ,  0�  |  0�  &  1[  &  1[  |  0�  |      C  , ,  0�  �  0�  F  1[  F  1[  �  0�  �      C  , ,  0�  �  0�  f  1[  f  1[  �  0�  �      C  , ,  0�   �  0�  �  1[  �  1[   �  0�   �      C  , ,  0�����  0�����  1[����  1[����  0�����      C  , ,  0����  0�����  1[����  1[���  0����      C  , ,  0����<  0�����  1[����  1[���<  0����<      C  , ,  0����\  0����  1[���  1[���\  0����\      C  , ,  0����|  0����&  1[���&  1[���|  0����|      C  , ,  0�����  0����F  1[���F  1[����  0�����      C  , ,  2  �  2  �  2�  �  2�  �  2  �      C  , ,  2    2  �  2�  �  2�    2        C  , ,  2  
<  2  
�  2�  
�  2�  
<  2  
<      C  , ,  2  \  2  	  2�  	  2�  \  2  \      C  , ,  2  |  2  &  2�  &  2�  |  2  |      C  , ,  2  �  2  F  2�  F  2�  �  2  �      C  , ,  2  �  2  f  2�  f  2�  �  2  �      C  , ,  2   �  2  �  2�  �  2�   �  2   �      C  , ,  2����  2����  2�����  2�����  2����      C  , ,  2���  2����  2�����  2����  2���      C  , ,  2���<  2����  2�����  2����<  2���<      ^   ,  .	����  .	  _  6�  _  6�����  .	����      A  , ,  *����b  *�  �  +�  �  +����b  *����b      A  , ,  +�  6  +�  �  9?  �  9?  6  +�  6      A  , ,  +����b  +����  9?���  9?���b  +����b      A  , ,  9?���b  9?  �  9�  �  9����b  9?���b      B  , ,  *�  �  *�  v  +�  v  +�  �  *�  �      B  , ,  9?  �  9?  v  9�  v  9�  �  9?  �      B  , ,  7A  �  7A  v  7�  v  7�  �  7A  �      B  , ,  9?  	�  9?  
n  9�  
n  9�  	�  9?  	�      B  , ,  9?  p  9?  	  9�  	  9�  p  9?  p      B  , ,  9?    9?  �  9�  �  9�    9?        B  , ,  9?  �  9?  r  9�  r  9�  �  9?  �      B  , ,  9?  t  9?    9�    9�  t  9?  t      B  , ,  9?     9?  �  9�  �  9�     9?         B  , ,  9?  l  9?    9�    9�  l  9?  l      B  , ,  9?  �  9?  j  9�  j  9�  �  9?  �      B  , ,  2�  6  2�  �  3m  �  3m  6  2�  6      B  , ,  2�  �  2�  �  3m  �  3m  �  2�  �      B  , ,  2�    2�  �  3m  �  3m    2�        B  , ,  2�  
<  2�  
�  3m  
�  3m  
<  2�  
<      B  , ,  2�  \  2�  	  3m  	  3m  \  2�  \      B  , ,  2�  |  2�  &  3m  &  3m  |  2�  |      B  , ,  2�  �  2�  F  3m  F  3m  �  2�  �      B  , ,  2�  �  2�  f  3m  f  3m  �  2�  �      B  , ,  7A  ,  7A  �  7�  �  7�  ,  7A  ,      B  , ,  4  6  4  �  4�  �  4�  6  4  6      B  , ,  4  �  4  �  4�  �  4�  �  4  �      B  , ,  4    4  �  4�  �  4�    4        B  , ,  4  
<  4  
�  4�  
�  4�  
<  4  
<      B  , ,  4  \  4  	  4�  	  4�  \  4  \      B  , ,  4  |  4  &  4�  &  4�  |  4  |      B  , ,  4  �  4  F  4�  F  4�  �  4  �      B  , ,  4  �  4  f  4�  f  4�  �  4  �      B  , ,  7A  l  7A    7�    7�  l  7A  l      B  , ,  5k  6  5k  �  6  �  6  6  5k  6      B  , ,  5k  �  5k  �  6  �  6  �  5k  �      B  , ,  5k    5k  �  6  �  6    5k        B  , ,  5k  
<  5k  
�  6  
�  6  
<  5k  
<      B  , ,  5k  \  5k  	  6  	  6  \  5k  \      B  , ,  5k  |  5k  &  6  &  6  |  5k  |      B  , ,  5k  �  5k  F  6  F  6  �  5k  �      B  , ,  5k  �  5k  f  6  f  6  �  5k  �      B  , ,  7A  �  7A  V  7�  V  7�  �  7A  �      B  , ,  6�  6  6�  �  7i  �  7i  6  6�  6      B  , ,  7A    7A  �  7�  �  7�    7A        B  , ,  7A  	L  7A  	�  7�  	�  7�  	L  7A  	L      B  , ,  7A  �  7A  6  7�  6  7�  �  7A  �      B  , ,  9?    9?  �  9�  �  9�    9?        B  , ,  -s  6  -s  �  .  �  .  6  -s  6      B  , ,  1o  6  1o  �  2  �  2  6  1o  6      B  , ,  .�  6  .�  �  /q  �  /q  6  .�  6      B  , ,  .�  �  .�  �  /q  �  /q  �  .�  �      B  , ,  .�    .�  �  /q  �  /q    .�        B  , ,  .�  
<  .�  
�  /q  
�  /q  
<  .�  
<      B  , ,  .�  \  .�  	  /q  	  /q  \  .�  \      B  , ,  .�  |  .�  &  /q  &  /q  |  .�  |      B  , ,  .�  �  .�  F  /q  F  /q  �  .�  �      B  , ,  .�  �  .�  f  /q  f  /q  �  .�  �      B  , ,  *�  �  *�  j  +�  j  +�  �  *�  �      B  , ,  *�  l  *�    +�    +�  l  *�  l      B  , ,  *�    *�  �  +�  �  +�    *�        B  , ,  *�  	�  *�  
n  +�  
n  +�  	�  *�  	�      B  , ,  *�  p  *�  	  +�  	  +�  p  *�  p      B  , ,  *�    *�  �  +�  �  +�    *�        B  , ,  *�  �  *�  r  +�  r  +�  �  *�  �      B  , ,  *�  t  *�    +�    +�  t  *�  t      B  , ,  0  6  0  �  0�  �  0�  6  0  6      B  , ,  0  �  0  �  0�  �  0�  �  0  �      B  , ,  0    0  �  0�  �  0�    0        B  , ,  0  
<  0  
�  0�  
�  0�  
<  0  
<      B  , ,  0  \  0  	  0�  	  0�  \  0  \      B  , ,  0  |  0  &  0�  &  0�  |  0  |      B  , ,  0  �  0  F  0�  F  0�  �  0  �      B  , ,  0  �  0  f  0�  f  0�  �  0  �      B  , ,  1o  �  1o  �  2  �  2  �  1o  �      B  , ,  1o    1o  �  2  �  2    1o        B  , ,  1o  
<  1o  
�  2  
�  2  
<  1o  
<      B  , ,  1o  \  1o  	  2  	  2  \  1o  \      B  , ,  1o  |  1o  &  2  &  2  |  1o  |      B  , ,  1o  �  1o  F  2  F  2  �  1o  �      B  , ,  1o  �  1o  f  2  f  2  �  1o  �      B  , ,  *�     *�  �  +�  �  +�     *�         B  , ,  1o���<  1o����  2����  2���<  1o���<      B  , ,  1o���\  1o���  2���  2���\  1o���\      B  , ,  1o���|  1o���&  2���&  2���|  1o���|      B  , ,  1o����  1o���F  2���F  2����  1o����      B  , ,  1o���b  1o���  2���  2���b  1o���b      B  , ,  0   �  0  �  0�  �  0�   �  0   �      B  , ,  *�   x  *�  "  +�  "  +�   x  *�   x      B  , ,  .�   �  .�  �  /q  �  /q   �  .�   �      B  , ,  0���\  0���  0����  0����\  0���\      B  , ,  0���|  0���&  0����&  0����|  0���|      B  , ,  0����  0���F  0����F  0�����  0����      B  , ,  0���b  0���  0����  0����b  0���b      B  , ,  *����|  *����&  +����&  +����|  *����|      B  , ,  *����(  *�����  +�����  +����(  *����(      B  , ,  *�����  *����~  +����~  +�����  *�����      B  , ,  *�����  *����*  +����*  +�����  *�����      B  , ,  *����,  *�����  +�����  +����,  *����,      B  , ,  *�����  *�����  +�����  +�����  *�����      B  , ,  -s���b  -s���  .���  .���b  -s���b      B  , ,  *����$  *�����  +�����  +����$  *����$      B  , ,  .�����  .�����  /q����  /q����  .�����      B  , ,  .����  .�����  /q����  /q���  .����      B  , ,  .����<  .�����  /q����  /q���<  .����<      B  , ,  .����\  .����  /q���  /q���\  .����\      B  , ,  .����|  .����&  /q���&  /q���|  .����|      B  , ,  .�����  .����F  /q���F  /q����  .�����      B  , ,  .����b  .����  /q���  /q���b  .����b      B  , ,  *�����  *����z  +����z  +�����  *�����      B  , ,  0����  0����  0�����  0�����  0����      B  , ,  0���  0����  0�����  0����  0���      B  , ,  0���<  0����  0�����  0����<  0���<      B  , ,  1o   �  1o  �  2  �  2   �  1o   �      B  , ,  1o����  1o����  2����  2����  1o����      B  , ,  1o���  1o����  2����  2���  1o���      B  , ,  5k���b  5k���  6���  6���b  5k���b      B  , ,  2����\  2����  3m���  3m���\  2����\      B  , ,  2����|  2����&  3m���&  3m���|  2����|      B  , ,  2�����  2����F  3m���F  3m����  2�����      B  , ,  2����b  2����  3m���  3m���b  2����b      B  , ,  7A���,  7A����  7�����  7����,  7A���,      B  , ,  2�   �  2�  �  3m  �  3m   �  2�   �      B  , ,  4   �  4  �  4�  �  4�   �  4   �      B  , ,  5k   �  5k  �  6  �  6   �  5k   �      B  , ,  9?   x  9?  "  9�  "  9�   x  9?   x      B  , ,  7A���l  7A���  7����  7����l  7A���l      B  , ,  9?����  9?����  9�����  9�����  9?����      B  , ,  6����b  6����  7i���  7i���b  6����b      B  , ,  7A���  7A����  7�����  7����  7A���      B  , ,  7A���L  7A����  7�����  7����L  7A���L      B  , ,  7A����  7A���6  7����6  7�����  7A����      B  , ,  9?���$  9?����  9�����  9����$  9?���$      B  , ,  9?����  9?���z  9����z  9�����  9?����      B  , ,  4����  4����  4�����  4�����  4����      B  , ,  4���  4����  4�����  4����  4���      B  , ,  4���<  4����  4�����  4����<  4���<      B  , ,  4���\  4���  4����  4����\  4���\      B  , ,  4���|  4���&  4����&  4����|  4���|      B  , ,  4����  4���F  4����F  4�����  4����      B  , ,  4���b  4���  4����  4����b  4���b      B  , ,  9?���|  9?���&  9����&  9����|  9?���|      B  , ,  9?���(  9?����  9�����  9����(  9?���(      B  , ,  9?����  9?���~  9����~  9�����  9?����      B  , ,  9?����  9?���*  9����*  9�����  9?����      B  , ,  9?���,  9?����  9�����  9����,  9?���,      B  , ,  7A����  7A   �  7�   �  7�����  7A����      B  , ,  2�����  2�����  3m����  3m����  2�����      B  , ,  2����  2�����  3m����  3m���  2����      B  , ,  2����<  2�����  3m����  3m���<  2����<      B  , ,  5k����  5k����  6����  6����  5k����      B  , ,  5k���  5k����  6����  6���  5k���      B  , ,  5k���<  5k����  6����  6���<  5k���<      B  , ,  5k���\  5k���  6���  6���\  5k���\      B  , ,  5k���|  5k���&  6���&  6���|  5k���|      B  , ,  5k����  5k���F  6���F  6����  5k����      @   ,  *?���  *?  �  :�  �  :����  *?���      A   ,  .����`  .�  �  6V  �  6V���`  .����`      ]  , ,  *v����  *v  ]  ,  ]  ,����  *v����      ]  , ,  ,  �  ,  ]  8�  ]  8�  �  ,  �      ]  , ,  ,����  ,���  8����  8�����  ,����      ]  , ,  8�����  8�  ]  :f  ]  :f����  8�����     �     0�     0 "sky130_fd_pr__nfet_01v8_P8PFL4    B   ,  �  �  �  �  (  �  (  �  �  �      B   ,���  ����  &  �  &  �  ����  �      B   ,  �    �  `  (  `  (    �        B   ,  �  6  �  �  (  �  (  6  �  6      B   ,���  p���    �    �  p���  p      B   ,���  P���  �  �  �  �  P���  P      B   ,  �  �  �     (     (  �  �  �      B   ,  �  �  �  @  (  @  (  �  �  �      B   ,���  0���  �  �  �  �  0���  0      B   ,���  	���  	�  �  	�  �  	���  	      B   ,  �  
�  �  �  (  �  (  
�  �  
�      B   ,  �  �  �  
   (  
   (  �  �  �      B   ,���  
����  �  �  �  �  
����  
�      B   ,���  ����  f  �  f  �  ����  �      B   ,  �  V  �  �  (  �  (  V  �  V      B   ,  �  v  �  �  (  �  (  v  �  v      B   ,���  ����  F  �  F  �  ����  �      B   ,���  ����  &  �  &  �  ����  �      B   ,  �    �  `  (  `  (    �        B   ,  �  6  �  �  (  �  (  6  �  6      B   ,���  p���    �    �  p���  p      B   ,���  P���  �  �  �  �  P���  P      B   ,  �  �  �     (     (  �  �  �      B   ,  �  �  �  @  (  @  (  �  �  �      B   ,���  0���  �  �  �  �  0���  0      B   ,���  ���  �  �  �  �  ���        B   ,  �  �  �     (     (  �  �  �      _   ,  �  "  �    <    <  "  �  "      C   ,���:���\���:  �����  ��������\���:���\      C   ,�������\�������  ,���  ,���\�������\      C   ,  .    .  `  �  `  �    .        C   ,  .  �  .     �     �  �  .  �      C   ,  .  
�  .  �  �  �  �  
�  .  
�      C   ,  .  V  .  �  �  �  �  V  .  V      C   ,  .    .  `  �  `  �    .        C   ,  .  �  .     �     �  �  .  �      C   ,����   �����  @  �  @  �   �����   �      C   ,����  v����     �     �  v����  v      C   ,����  V����     �     �  V����  V      C   ,����  6����  �  �  �  �  6����  6      C   ,����  ����  �  �  �  �  ����        C   ,����  	�����  
�  �  
�  �  	�����  	�      C   ,����  �����  �  �  �  �  �����  �      C   ,����  �����  `  �  `  �  �����  �      C   ,����  �����  @  �  @  �  �����  �      C   ,����  v����     �     �  v����  v      C   ,����  V����     �     �  V����  V      C   ,����  6����  �  �  �  �  6����  6      C   ,����  ����  �  �  �  �  ����        C   ,����  �����  �  �  �  �  �����  �      C   ,  .  6  .  �  �  �  �  6  .  6      C   ,  .  �  .  @  �  @  �  �  .  �      C   ,  .  �  .  
   �  
   �  �  .  �      C   ,  .  v  .  �  �  �  �  v  .  v      C   ,  .  6  .  �  �  �  �  6  .  6      C   ,  .  �  .  @  �  @  �  �  .  �      C   ,  .  �  .     �     �  �  .  �      C   ,����  0����  �  ,  �  ,  0����  0      C   ,  ,���\  ,  �  �  �  ����\  ,���\      C   ,  .  �  .  �  �  �  �  �  .  �      D   ,    *    L  �  L  �  *    *      D   ,    �      �    �  �    �      D   ,    
�    �  �  �  �  
�    
�      D   ,    j    �  �  �  �  j    j      D   ,    *    L  �  L  �  *    *      D   ,    �      �    �  �    �      D   ,���u   x���u  ^  E  ^  E   x���u   x      D   ,���u  X���u  >  E  >  E  X���u  X      D   ,����  8����    p    p  8����  8      D   ,���u  ���u  �  E  �  E  ���u        D   ,����  �����  �  p  �  p  �����  �      D   ,���u  	����u  
�  E  
�  E  	����u  	�      D   ,����  �����  �  p  �  p  �����  �      D   ,���u  ����u  ~  E  ~  E  ����u  �      D   ,����  x����  ^  p  ^  p  x����  x      D   ,���u  X���u  >  E  >  E  X���u  X      D   ,����  8����    p    p  8����  8      D   ,���u  ���u  �  E  �  E  ���u        D   ,����  �����  �  p  �  p  �����  �      D   ,����  �����  �  p  �  p  �����  �      D   ,    J    l  �  l  �  J    J      D   ,    
    ,  �  ,  �  
    
      D   ,    �    	�  �  	�  �  �    �      D   ,    �    �  �  �  �  �    �      D   ,    J    l  �  l  �  J    J      D   ,    
    ,  �  ,  �  
    
      D   ,    �    �  �  �  �  �    �      D   ,    J    �  x  �  x  J    J      C  , ,  .  f  .    �    �  f  .  f      C  , ,  .  &  .  �  �  �  �  &  .  &      C  , ,  .  
�  .  �  �  �  �  
�  .  
�      C  , ,  .  �  .  P  �  P  �  �  .  �      C  , ,  .  f  .    �    �  f  .  f      C  , ,  .  &  .  �  �  �  �  &  .  &      C  , ,���c   ����c  @���  @���   ����c   �      C  , ,���c  v���c   ���   ���  v���c  v      C  , ,���c  V���c   ���   ���  V���c  V      C  , ,���c  6���c  ����  ����  6���c  6      C  , ,���c  ���c  ����  ����  ���c        C  , ,���c  	����c  
����  
����  	����c  	�      C  , ,���c  ����c  ����  ����  ����c  �      C  , ,���c  ����c  `���  `���  ����c  �      C  , ,���c  ����c  @���  @���  ����c  �      C  , ,���c  v���c   ���   ���  v���c  v      C  , ,���c  V���c   ���   ���  V���c  V      C  , ,���c  6���c  ����  ����  6���c  6      C  , ,���c  ���c  ����  ����  ���c        C  , ,���c  ����c  ����  ����  ����c  �      C  , ,����   �����  @���u  @���u   �����   �      C  , ,����  v����   ���u   ���u  v����  v      C  , ,����  V����   ���u   ���u  V����  V      C  , ,����  6����  ����u  ����u  6����  6      C  , ,����  ����  ����u  ����u  ����        C  , ,����  	�����  
����u  
����u  	�����  	�      C  , ,����  �����  ����u  ����u  �����  �      C  , ,����  �����  `���u  `���u  �����  �      C  , ,����  �����  @���u  @���u  �����  �      C  , ,����  v����   ���u   ���u  v����  v      C  , ,����  V����   ���u   ���u  V����  V      C  , ,����  6����  ����u  ����u  6����  6      C  , ,����  ����  ����u  ����u  ����        C  , ,����  �����  ����u  ����u  �����  �      C  , ,���3   ����3  @����  @����   ����3   �      C  , ,���3  v���3   ����   ����  v���3  v      C  , ,���3  V���3   ����   ����  V���3  V      C  , ,���3  6���3  �����  �����  6���3  6      C  , ,���3  ���3  �����  �����  ���3        C  , ,���3  	����3  
�����  
�����  	����3  	�      C  , ,���3  ����3  �����  �����  ����3  �      C  , ,���3  ����3  `����  `����  ����3  �      C  , ,���3  ����3  @����  @����  ����3  �      C  , ,���3  v���3   ����   ����  v���3  v      C  , ,���3  V���3   ����   ����  V���3  V      C  , ,���3  6���3  �����  �����  6���3  6      C  , ,���3  ���3  �����  �����  ���3        C  , ,���3  ����3  �����  �����  ����3  �      C  , ,   �  V   �     E     E  V   �  V      C  , ,   �     �  �  E  �  E     �        C  , ,   �  �   �  �  E  �  E  �   �  �      C  , ,   �  �   �  @  E  @  E  �   �  �      C  , ,   �  V   �     E     E  V   �  V      C  , ,   �     �  �  E  �  E     �        C  , ,   �  �   �  �  E  �  E  �   �  �      C  , ,    V       �     �  V    V      C  , ,        �  �  �  �            C  , ,    �    �  �  �  �  �    �      C  , ,    �    @  �  @  �  �    �      C  , ,    V       �     �  V    V      C  , ,        �  �  �  �            C  , ,    �    �  �  �  �  �    �      C  , ,  .  �  .  0  �  0  �  �  .  �      C  , ,  .  F  .  �  �  �  �  F  .  F      C  , ,  .  	  .  	�  �  	�  �  	  .  	      C  , ,  .  �  .  p  �  p  �  �  .  �      C  , ,  .  �  .  0  �  0  �  �  .  �      C  , ,  .  F  .  �  �  �  �  F  .  F      C  , ,  .    .  �  �  �  �    .        ^   ,������������  W���a  W���a������������      ^   ,���a�������a����  �����  ��������a����      ^   ,���a  ����a  W  �  W  �  ����a  �      ^   ,  �����  �  W  S  W  S����  �����      A  , ,���:���\���:  �����  ��������\���:���\      A  , ,�������\�������  ,���  ,���\�������\      A  , ,����  0����  �  ,  �  ,  0����  0      A  , ,  ,���\  ,  �  �  �  ����\  ,���\      B  , ,  ,  �  ,  p  �  p  �  �  ,  �      B  , ,  .  �  .  p  �  p  �  �  .  �      B  , ,���:  ����:  p����  p����  ����:  �      B  , ,  .    .  �  �  �  �    .        B  , ,  �  0  �  �  �  �  �  0  �  0      B  , ,  .  �  .  0  �  0  �  �  .  �      B  , ,  1  �  1  �  �  �  �  �  1  �      B  , ,  ,    ,  �  �  �  �    ,        B  , ,  ,  n  ,    �    �  n  ,  n      B  , ,  ,  �  ,  l  �  l  �  �  ,  �      B  , ,  �  �  �  `  /  `  /  �  �  �      B  , ,  �  �  �  @  /  @  /  �  �  �      B  , ,  �  v  �     /     /  v  �  v      B  , ,  �  V  �     /     /  V  �  V      B  , ,  �  6  �  �  /  �  /  6  �  6      B  , ,  �    �  �  /  �  /    �        B  , ,  �  �  �  �  /  �  /  �  �  �      B  , ,  �  0  �  �  /  �  /  0  �  0      B  , ,  ,    ,  �  �  �  �    ,        B  , ,  .  �  .  P  �  P  �  �  .  �      B  , ,  .  f  .    �    �  f  .  f      B  , ,  .  &  .  �  �  �  �  &  .  &      B  , ,  1  0  1  �  �  �  �  0  1  0      B  , ,����  �����  `   �  `   �  �����  �      B  , ,����  �����  @   �  @   �  �����  �      B  , ,����  v����      �      �  v����  v      B  , ,����  V����      �      �  V����  V      B  , ,����  6����  �   �  �   �  6����  6      B  , ,����  ����  �   �  �   �  ����        B  , ,����  �����  �   �  �   �  �����  �      B  , ,����  0����  �   �  �   �  0����  0      B  , ,  .  F  .  �  �  �  �  F  .  F      B  , ,  ,  j  ,    �    �  j  ,  j      B  , ,  ,  �  ,  h  �  h  �  �  ,  �      B  , ,  ,    ,  �  �  �  �    ,        B  , ,  ,  f  ,    �    �  f  ,  f      B  , ,  ,  �  ,  d  �  d  �  �  ,  �      B  , ,  1  �  1  `  �  `  �  �  1  �      B  , ,  1  �  1  @  �  @  �  �  1  �      B  , ,  1  v  1     �     �  v  1  v      B  , ,  1  V  1     �     �  V  1  V      B  , ,  1  6  1  �  �  �  �  6  1  6      B  , ,  1    1  �  �  �  �    1        B  , ,����  V����   ���3   ���3  V����  V      B  , ,����  6����  ����3  ����3  6����  6      B  , ,����  ����  ����3  ����3  ����        B  , ,����  �����  ����3  ����3  �����  �      B  , ,����  0����  ����3  ����3  0����  0      B  , ,���:  ����:  l����  l����  ����:  �      B  , ,���:  ���:  �����  �����  ���:        B  , ,���:  j���:  ����  ����  j���:  j      B  , ,���:  ����:  h����  h����  ����:  �      B  , ,���:  ���:  �����  �����  ���:        B  , ,���:  f���:  ����  ����  f���:  f      B  , ,���:  ����:  d����  d����  ����:  �      B  , ,����  0����  ����7  ����7  0����  0      B  , ,���5  ����5  `����  `����  ����5  �      B  , ,����  �����  `����  `����  �����  �      B  , ,����  �����  @����  @����  �����  �      B  , ,����  v����   ����   ����  v����  v      B  , ,����  V����   ����   ����  V����  V      B  , ,����  6����  �����  �����  6����  6      B  , ,����  ����  �����  �����  ����        B  , ,����  �����  �����  �����  �����  �      B  , ,����  0����  �����  �����  0����  0      B  , ,���:  ���:  �����  �����  ���:        B  , ,���5  ����5  @����  @����  ����5  �      B  , ,���5  v���5   ����   ����  v���5  v      B  , ,���5  V���5   ����   ����  V���5  V      B  , ,���5  6���5  �����  �����  6���5  6      B  , ,���5  ���5  �����  �����  ���5        B  , ,���5  ����5  �����  �����  ����5  �      B  , ,���5  0���5  �����  �����  0���5  0      B  , ,���:  n���:  ����  ����  n���:  n      B  , ,����  �����  `���3  `���3  �����  �      B  , ,����  �����  @���3  @���3  �����  �      B  , ,����  v����   ���3   ���3  v����  v      B  , ,���:  z���:  $����  $����  z���:  z      B  , ,�������\����������7������7���\�������\      B  , ,���:  ����:  x����  x����  ����:  �      B  , ,���5���\���5�����������������\���5���\      B  , ,���5   ����5  @����  @����   ����5   �      B  , ,���5  v���5   ����   ����  v���5  v      B  , ,���5  V���5   ����   ����  V���5  V      B  , ,���5  6���5  �����  �����  6���5  6      B  , ,���5  ���5  �����  �����  ���5        B  , ,���5  	����5  
�����  
�����  	����5  	�      B  , ,�������\���������������������\�������\      B  , ,����   �����  @����  @����   �����   �      B  , ,����  v����   ����   ����  v����  v      B  , ,����  V����   ����   ����  V����  V      B  , ,����  6����  �����  �����  6����  6      B  , ,����  ����  �����  �����  ����        B  , ,����  	�����  
�����  
�����  	�����  	�      B  , ,���:  "���:  �����  �����  "���:  "      B  , ,���:  v���:   ����   ����  v���:  v      B  , ,�������\����������3������3���\�������\      B  , ,����   �����  @���3  @���3   �����   �      B  , ,����  v����   ���3   ���3  v����  v      B  , ,����  V����   ���3   ���3  V����  V      B  , ,����  �����  ����3  ����3  �����  �      B  , ,���:  r���:  ����  ����  r���:  r      B  , ,����  �����  �����  �����  �����  �      B  , ,���5  ����5  �����  �����  ����5  �      B  , ,����  6����  ����3  ����3  6����  6      B  , ,����  ����  ����3  ����3  ����        B  , ,����  	�����  
����3  
����3  	�����  	�      B  , ,���:  ����:  	t����  	t����  ����:  �      B  , ,���:  
���:  
�����  
�����  
���:  
      B  , ,���:   ����:  |����  |����   ����:   �      B  , ,���:  &���:  �����  �����  &���:  &      B  , ,  ,  �  ,  	t  �  	t  �  �  ,  �      B  , ,  ,  
  ,  
�  �  
�  �  
  ,  
      B  , ,  ,   �  ,  |  �  |  �   �  ,   �      B  , ,  ,  &  ,  �  �  �  �  &  ,  &      B  , ,  ,  z  ,  $  �  $  �  z  ,  z      B  , ,  ,  �  ,  x  �  x  �  �  ,  �      B  , ,  ,  "  ,  �  �  �  �  "  ,  "      B  , ,  .  f  .    �    �  f  .  f      B  , ,  .  &  .  �  �  �  �  &  .  &      B  , ,  1���\  1���  ����  ����\  1���\      B  , ,  1   �  1  @  �  @  �   �  1   �      B  , ,  1  v  1     �     �  v  1  v      B  , ,  1  V  1     �     �  V  1  V      B  , ,  1  6  1  �  �  �  �  6  1  6      B  , ,  1    1  �  �  �  �    1        B  , ,  1  	�  1  
�  �  
�  �  	�  1  	�      B  , ,  .  
�  .  �  �  �  �  
�  .  
�      B  , ,  ����\  ����  /���  /���\  ����\      B  , ,  �   �  �  @  /  @  /   �  �   �      B  , ,  �  v  �     /     /  v  �  v      B  , ,  �  V  �     /     /  V  �  V      B  , ,  �  6  �  �  /  �  /  6  �  6      B  , ,  �    �  �  /  �  /    �        B  , ,  �  	�  �  
�  /  
�  /  	�  �  	�      B  , ,  ,  v  ,     �     �  v  ,  v      B  , ,  ����\  ����  ����  ����\  ����\      B  , ,  .  �  .  0  �  0  �  �  .  �      B  , ,  .  F  .  �  �  �  �  F  .  F      B  , ,  .  	  .  	�  �  	�  �  	  .  	      B  , ,  �  �  �  �  /  �  /  �  �  �      B  , ,����  �����  �   �  �   �  �����  �      B  , ,  ,  r  ,    �    �  r  ,  r      B  , ,�������\�������   ����   ����\�������\      B  , ,����   �����  @   �  @   �   �����   �      B  , ,����  v����      �      �  v����  v      B  , ,����  V����      �      �  V����  V      B  , ,����  6����  �   �  �   �  6����  6      B  , ,����  ����  �   �  �   �  ����        B  , ,����  	�����  
�   �  
�   �  	�����  	�      B  , ,  1  �  1  �  �  �  �  �  1  �      A   ,����   Z����  �  p  �  p   Z����   Z      ]  , ,���#�������#  Y  �  Y  ��������#����     �     0�     0 "sky130_fd_pr__pfet_01v8_VCXY4M 
  via_new     B�       ����  �      B   ,  ����Q  �  >  ;  >  ;���Q  ����Q      B   ,  ����Q  �  >  [  >  [���Q  ����Q      B   ,  ����Q  �  >  {  >  {���Q  ����Q      B   ,  ���Q    >  �  >  ����Q  ���Q      B   ,  %���Q  %  >  �  >  ����Q  %���Q      B   ,  E���Q  E  >  �  >  ����Q  E���Q      B   ,  	e���Q  	e  >  	�  >  	����Q  	e���Q      B   ,  ����Q  �  >    >  ���Q  ����Q      B   ,  ����Q  �  >  ;  >  ;���Q  ����Q      B   ,  ����Q  �  >  [  >  [���Q  ����Q      B   ,  ����Q  �  >  {  >  {���Q  ����Q      B   ,   ���Q     >   �  >   ����Q   ���Q      B   ,���%���Q���%  >����  >�������Q���%���Q      B   ,����  >����  �  �  �  �  >����  >      B   ,  �  �  �  u  ;  u  ;  �  �  �      B   ,  �  �  �  u  [  u  [  �  �  �      B   ,  �  �  �  u  {  u  {  �  �  �      B   ,    �    u  �  u  �  �    �      B   ,  %  �  %  u  �  u  �  �  %  �      B   ,  E  �  E  u  �  u  �  �  E  �      B   ,  	e  �  	e  u  	�  u  	�  �  	e  �      B   ,  �  �  �  u    u    �  �  �      B   ,  �  �  �  u  ;  u  ;  �  �  �      B   ,  �  �  �  u  [  u  [  �  �  �      B   ,  �  �  �  u  {  u  {  �  �  �      B   ,     �     u   �  u   �  �     �      B   ,���%  ����%  u����  u����  ����%  �      C   ,�������@��������  o����  o���@�������@      C   ,  �����  �  �  5  �  5����  �����      C   ,  �����  �  �  U  �  U����  �����      C   ,  �����  �  �  u  �  u����  �����      C   ,  �����  �  �  �  �  �����  �����      C   ,  ����    �  �  �  �����  ����      C   ,  +����  +  �  �  �  �����  +����      C   ,  
K����  
K  �  
�  �  
�����  
K����      C   ,  k����  k  �  	  �  	����  k����      C   ,  �����  �  �  5  �  5����  �����      C   ,  �����  �  �  U  �  U����  �����      C   ,  �����  �  �  u  �  u����  �����      C   ,   �����   �  �  �  �  �����   �����      C   ,����������  �����  ����������������      C   ,���+�������+  �����  ������������+����      C   ,������������  �����  �����������������      C   ,  �����  �  �  o  �  o����  �����      C   ,����  �����  �  o  �  o  �����  �      C   ,  �    �    5    5    �        C   ,  �    �    U    U    �        C   ,  �    �    u    u    �        C   ,  �    �    �    �    �        C   ,          �    �            C   ,  +    +    �    �    +        C   ,  
K    
K    
�    
�    
K        C   ,  k    k    	    	    k        C   ,  �    �    5    5    �        C   ,  �    �    U    U    �        C   ,  �    �    u    u    �        C   ,   �     �    �    �     �        C   ,���  ���  ����  ����  ���        C   ,���+  ���+  ����  ����  ���+        D   ,  m����  m  �  S  �  S����  m����      D   ,  �����  �  �  s  �  s����  �����      D   ,  �����  �  �  �  �  �����  �����      D   ,  �����  �  �  �  �  �����  �����      D   ,  �����  �  �  �  �  �����  �����      D   ,  ����    �  �  �  �����  ����      D   ,  
-����  
-  �    �  ����  
-����      D   ,  M����  M  �  	3  �  	3����  M����      D   ,  m����  m  �  S  �  S����  m����      D   ,  �����  �  �  s  �  s����  �����      D   ,  �����  �  �  �  �  �����  �����      D   ,   �����   �  �  �  �  �����   �����      D   ,������������  �����  �����������������      D   ,����������  �����  ����������������      D   ,  m  #  m  �  S  �  S  #  m  #      D   ,  �  #  �  �  s  �  s  #  �  #      D   ,  �  #  �  �  �  �  �  #  �  #      D   ,  �  #  �  �  �  �  �  #  �  #      D   ,  �  #  �  �  �  �  �  #  �  #      D   ,    #    �  �  �  �  #    #      D   ,  
-  #  
-  �    �    #  
-  #      D   ,  M  #  M  �  	3  �  	3  #  M  #      D   ,  m  #  m  �  S  �  S  #  m  #      D   ,  �  #  �  �  s  �  s  #  �  #      D   ,  �  #  �  �  �  �  �  #  �  #      D   ,   �  #   �  �  �  �  �  #   �  #      D   ,����  #����  �����  �����  #����  #      D   ,���  #���  �����  �����  #���  #      D   ,  s����  s  �  m  �  m����  s����      D   ,  s  #  s  �  m  �  m  #  s  #      D   ,������������  �����  �����������������      D   ,����  #����  �����  �����  #����  #      D   ,   �  �   �  #  �  #  �  �   �  �      D   ,  �  �  �  #  s  #  s  �  �  �      D   ,  M  �  M  #  	3  #  	3  �  M  �      D   ,    �    #  �  #  �  �    �      D   ,  �  �  �  #  �  #  �  �  �  �      D   ,  �  �  �  #  s  #  s  �  �  �      D   ,   �  >   �  �  s  �  s  >   �  >      D   ,����  �����  -����  -����  �����  �      D   ,  �  �  �  -  �  -  �  �  �  �      D   ,  m  �  m  -  S  -  S  �  m  �      D   ,  
-  �  
-  -    -    �  
-  �      D   ,  �  �  �  -  �  -  �  �  �  �      D   ,  �  �  �  -  �  -  �  �  �  �      D   ,����  -����  ;  �  ;  �  -����  -      D   ,����������������������������������������      D   ,  �����  �����  �����  �����  �����      D   ,  m����  m����  S����  S����  m����      D   ,  
-����  
-����  ����  ����  
-����      D   ,  �����  �����  �����  �����  �����      D   ,  �����  �����  �����  �����  �����      D   ,����������������  �����  �������������      D   ,����  f����  `����  `����  f����  f      C  , ,  
K  �  
K  0  
�  0  
�  �  
K  �      C  , ,  �  �  �  �  5  �  5  �  �  �      C  , ,  �  �  �  �  U  �  U  �  �  �      C  , ,    N    �  �  �  �  N    N      C  , ,  +  N  +  �  �  �  �  N  +  N      C  , ,  
K  N  
K  �  
�  �  
�  N  
K  N      C  , ,  �  �  �  0  5  0  5  �  �  �      C  , ,  �  �  �  0  U  0  U  �  �  �      C  , ,  �  �  �  0  u  0  u  �  �  �      C  , ,  �  �  �  0  �  0  �  �  �  �      C  , ,    �    0  �  0  �  �    �      C  , ,  +  �  +  0  �  0  �  �  +  �      C  , ,    �    	`  �  	`  �  �    �      C  , ,  +  �  +  	`  �  	`  �  �  +  �      C  , ,  
K  �  
K  	`  
�  	`  
�  �  
K  �      C  , ,  �  �  �  �  u  �  u  �  �  �      C  , ,  �  �  �  �  �  �  �  �  �  �      C  , ,    �    �  �  �  �  �    �      C  , ,  +  �  +  �  �  �  �  �  +  �      C  , ,  
K  �  
K  �  
�  �  
�  �  
K  �      C  , ,  �  �  �  	`  5  	`  5  �  �  �      C  , ,  �  �  �  	`  U  	`  U  �  �  �      C  , ,  �  �  �  	`  u  	`  u  �  �  �      C  , ,  �  �  �  	`  �  	`  �  �  �  �      C  , ,  �  
  �  
�  5  
�  5  
  �  
      C  , ,  �  
  �  
�  U  
�  U  
  �  
      C  , ,  �  
  �  
�  u  
�  u  
  �  
      C  , ,  �  
  �  
�  �  
�  �  
  �  
      C  , ,    
    
�  �  
�  �  
    
      C  , ,  +  
  +  
�  �  
�  �  
  +  
      C  , ,  
K  
  
K  
�  
�  
�  
�  
  
K  
      C  , ,  �  N  �  �  5  �  5  N  �  N      C  , ,  �  N  �  �  U  �  U  N  �  N      C  , ,  �  N  �  �  u  �  u  N  �  N      C  , ,  �  N  �  �  �  �  �  N  �  N      C  , ,  k  �  k  0  	  0  	  �  k  �      C  , ,  �  �  �  0  5  0  5  �  �  �      C  , ,  �  �  �  0  U  0  U  �  �  �      C  , ,  �  �  �  0  u  0  u  �  �  �      C  , ,   �  �   �  0  �  0  �  �   �  �      C  , ,���  ����  0����  0����  ����  �      C  , ,���+  ����+  0����  0����  ����+  �      C  , ,  k  
  k  
�  	  
�  	  
  k  
      C  , ,  �  
  �  
�  5  
�  5  
  �  
      C  , ,  �  
  �  
�  U  
�  U  
  �  
      C  , ,  �  
  �  
�  u  
�  u  
  �  
      C  , ,   �  
   �  
�  �  
�  �  
   �  
      C  , ,���  
���  
�����  
�����  
���  
      C  , ,���+  
���+  
�����  
�����  
���+  
      C  , ,  k  �  k  	`  	  	`  	  �  k  �      C  , ,  �  �  �  	`  5  	`  5  �  �  �      C  , ,  �  �  �  	`  U  	`  U  �  �  �      C  , ,  �  �  �  	`  u  	`  u  �  �  �      C  , ,   �  �   �  	`  �  	`  �  �   �  �      C  , ,���  ����  	`����  	`����  ����  �      C  , ,���+  ����+  	`����  	`����  ����+  �      C  , ,  k  N  k  �  	  �  	  N  k  N      C  , ,  �  N  �  �  5  �  5  N  �  N      C  , ,  �  N  �  �  U  �  U  N  �  N      C  , ,  �  N  �  �  u  �  u  N  �  N      C  , ,   �  N   �  �  �  �  �  N   �  N      C  , ,���  N���  �����  �����  N���  N      C  , ,���+  N���+  �����  �����  N���+  N      C  , ,  k  �  k  �  	  �  	  �  k  �      C  , ,  �  �  �  �  5  �  5  �  �  �      C  , ,  �  �  �  �  U  �  U  �  �  �      C  , ,  �  �  �  �  u  �  u  �  �  �      C  , ,   �  �   �  �  �  �  �  �   �  �      C  , ,���  ����  �����  �����  ����  �      C  , ,���+  ����+  �����  �����  ����+  �      C  , ,  k����  k���@  	���@  	����  k����      C  , ,  �����  ����@  5���@  5����  �����      C  , ,  �����  ����@  U���@  U����  �����      C  , ,  �����  ����@  u���@  u����  �����      C  , ,   �����   ����@  ����@  �����   �����      C  , ,�������������@�������@���������������      C  , ,���+�������+���@�������@�����������+����      C  , ,  k����  k����  	����  	����  k����      C  , ,  �����  �����  5����  5����  �����      C  , ,  �����  �����  U����  U����  �����      C  , ,  �����  �����  u����  u����  �����      C  , ,   �����   �����  �����  �����   �����      C  , ,�������������������������������������      C  , ,���+�������+�����������������������+����      C  , ,  k���f  k���  	���  	���f  k���f      C  , ,  ����f  ����  5���  5���f  ����f      C  , ,  ����f  ����  U���  U���f  ����f      C  , ,  ����f  ����  u���  u���f  ����f      C  , ,   ����f   ����  ����  ����f   ����f      C  , ,������f��������������������f������f      C  , ,���+���f���+�����������������f���+���f      C  , ,  k����  k   x  	   x  	����  k����      C  , ,  �����  �   x  5   x  5����  �����      C  , ,  �����  �   x  U   x  U����  �����      C  , ,  �����  �   x  u   x  u����  �����      C  , ,   �����   �   x  �   x  �����   �����      C  , ,����������   x����   x���������������      C  , ,���+�������+   x����   x�����������+����      C  , ,  k  6  k  �  	  �  	  6  k  6      C  , ,  �  6  �  �  5  �  5  6  �  6      C  , ,  �  6  �  �  U  �  U  6  �  6      C  , ,  �  6  �  �  u  �  u  6  �  6      C  , ,   �  6   �  �  �  �  �  6   �  6      C  , ,���  6���  �����  �����  6���  6      C  , ,���+  6���+  �����  �����  6���+  6      C  , ,  �����  �����  5����  5����  �����      C  , ,  �����  �����  U����  U����  �����      C  , ,  �����  �����  u����  u����  �����      C  , ,  �����  �����  �����  �����  �����      C  , ,  ����  ����  �����  �����  ����      C  , ,  +����  +����  �����  �����  +����      C  , ,  
K����  
K����  
�����  
�����  
K����      C  , ,  �����  �   x  5   x  5����  �����      C  , ,  �����  �   x  U   x  U����  �����      C  , ,  �����  �   x  u   x  u����  �����      C  , ,  �����  �   x  �   x  �����  �����      C  , ,  ����     x  �   x  �����  ����      C  , ,  +����  +   x  �   x  �����  +����      C  , ,  
K����  
K   x  
�   x  
�����  
K����      C  , ,  �����  ����@  5���@  5����  �����      C  , ,  �����  ����@  U���@  U����  �����      C  , ,  �����  ����@  u���@  u����  �����      C  , ,  �����  ����@  ����@  �����  �����      C  , ,  ����  ���@  ����@  �����  ����      C  , ,  +����  +���@  ����@  �����  +����      C  , ,  
K����  
K���@  
����@  
�����  
K����      C  , ,  �  6  �  �  5  �  5  6  �  6      C  , ,  �  6  �  �  U  �  U  6  �  6      C  , ,  �  6  �  �  u  �  u  6  �  6      C  , ,  �  6  �  �  �  �  �  6  �  6      C  , ,    6    �  �  �  �  6    6      C  , ,  +  6  +  �  �  �  �  6  +  6      C  , ,  
K  6  
K  �  
�  �  
�  6  
K  6      C  , ,  ����f  ����  5���  5���f  ����f      C  , ,  ����f  ����  U���  U���f  ����f      C  , ,  ����f  ����  u���  u���f  ����f      C  , ,  ����f  ����  ����  ����f  ����f      C  , ,  ���f  ���  ����  ����f  ���f      C  , ,  +���f  +���  ����  ����f  +���f      C  , ,  
K���f  
K���  
����  
����f  
K���f      ^   ,���r���V���r     �     ����V���r���V      ^   ,���r  ����r  p  �  p  �  ����r  �      A  , ,����  �����  �  o  �  o  �����  �      A  , ,  �  :  �  �  o  �  o  :  �  :      A  , ,����  :����  �����  �����  :����  :      A  , ,�������@��������  o����  o���@�������@      A  , ,  �����  �  �  o  �  o����  �����      A  , ,������������  �����  �����������������      B  , ,���+  ����+  8����  8����  ����+  �      B  , ,  	[���@  	[����  
����  
���@  	[���@      B  , ,  	[  �  	[  �  
  �  
  �  	[  �      B  , ,  +  d  +    �    �  d  +  d      B  , ,  �    �  �  o  �  o    �        B  , ,  �    �  �  5  �  5    �        B  , ,  �    �  �  U  �  U    �        B  , ,  �    �  �  u  �  u    �        B  , ,  �    �  �  �  �  �    �        B  , ,        �  �  �  �            B  , ,  +    +  �  �  �  �    +        B  , ,  �  
�  �  ^  �  ^  �  
�  �  
�      B  , ,    
�    ^  �  ^  �  
�    
�      B  , ,  +  
�  +  ^  �  ^  �  
�  +  
�      B  , ,  
K  
�  
K  ^  
�  ^  
�  
�  
K  
�      B  , ,  �  \  �    o    o  \  �  \      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �    �  �  o  �  o    �        B  , ,  �    �  �  5  �  5    �        B  , ,  �    �  �  U  �  U    �        B  , ,  �    �  �  u  �  u    �        B  , ,  �    �  �  �  �  �    �        B  , ,        �  �  �  �            B  , ,  +    +  �  �  �  �    +        B  , ,  
K    
K  �  
�  �  
�    
K        B  , ,  �  �  �  �  Q  �  Q  �  �  �      B  , ,  S  �  S  �  �  �  �  �  S  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  �  �  �  U  �  U  �  �  �      B  , ,  W  �  W  �    �    �  W  �      B  , ,    �    �  �  �  �  �    �      B  , ,  
�  �  
�  �  Y  �  Y  �  
�  �      B  , ,  O  �  O  �  �  �  �  �  O  �      B  , ,  �  
�  �  ^  o  ^  o  
�  �  
�      B  , ,  �  
�  �  ^  5  ^  5  
�  �  
�      B  , ,  �  
�  �  ^  U  ^  U  
�  �  
�      B  , ,  �  
�  �  ^  u  ^  u  
�  �  
�      B  , ,  
K  d  
K    
�    
�  d  
K  d      B  , ,  
K  �  
K  b  
�  b  
�  �  
K  �      B  , ,  
K    
K  �  
�  �  
�    
K        B  , ,  �  �  �  b  o  b  o  �  �  �      B  , ,  �  �  �  b  5  b  5  �  �  �      B  , ,  �  �  �  b  U  b  U  �  �  �      B  , ,  �  �  �  b  u  b  u  �  �  �      B  , ,  �  �  �  b  �  b  �  �  �  �      B  , ,    �    b  �  b  �  �    �      B  , ,  �  	`  �  

  o  

  o  	`  �  	`      B  , ,  �  	`  �  

  5  

  5  	`  �  	`      B  , ,  �  	`  �  

  U  

  U  	`  �  	`      B  , ,  �  	`  �  

  u  

  u  	`  �  	`      B  , ,  �  	`  �  

  �  

  �  	`  �  	`      B  , ,    	`    

  �  

  �  	`    	`      B  , ,  +  	`  +  

  �  

  �  	`  +  	`      B  , ,  
K  	`  
K  

  
�  

  
�  	`  
K  	`      B  , ,  +  �  +  b  �  b  �  �  +  �      B  , ,  �  d  �    o    o  d  �  d      B  , ,  �  d  �    5    5  d  �  d      B  , ,  �  d  �    U    U  d  �  d      B  , ,  �  d  �    u    u  d  �  d      B  , ,  �  d  �    �    �  d  �  d      B  , ,    d      �    �  d    d      B  , ,  k  	`  k  

  	  

  	  	`  k  	`      B  , ,���g  ����g  ����  ����  ����g  �      B  , ,����  \����  ����  ����  \����  \      B  , ,  k    k  �  	  �  	    k        B  , ,  �    �  �  5  �  5    �        B  , ,  �    �  �  U  �  U    �        B  , ,  �    �  �  u  �  u    �        B  , ,   �     �  �  �  �  �     �        B  , ,���  ���  �����  �����  ���        B  , ,���+  ���+  �����  �����  ���+        B  , ,����  ����  �����  �����  ����        B  , ,  k  
�  k  ^  	  ^  	  
�  k  
�      B  , ,  �  
�  �  ^  5  ^  5  
�  �  
�      B  , ,  �  
�  �  ^  U  ^  U  
�  �  
�      B  , ,  �  
�  �  ^  u  ^  u  
�  �  
�      B  , ,   �  
�   �  ^  �  ^  �  
�   �  
�      B  , ,���  
����  ^����  ^����  
����  
�      B  , ,���+  
����+  ^����  ^����  
����+  
�      B  , ,����  
�����  ^����  ^����  
�����  
�      B  , ,    �    �  �  �  �  �    �      B  , ,  �  �  �  �  ]  �  ]  �  �  �      B  , ,  _  �  _  �  	  �  	  �  _  �      B  , ,    �    �  �  �  �  �    �      B  , ,  �  �  �  �  a  �  a  �  �  �      B  , ,  c  �  c  �    �    �  c  �      B  , ,     �     �   �  �   �  �     �      B  , ,����  �����  ����e  ����e  �����  �      B  , ,  �  	`  �  

  5  

  5  	`  �  	`      B  , ,  �  	`  �  

  U  

  U  	`  �  	`      B  , ,  �  	`  �  

  u  

  u  	`  �  	`      B  , ,   �  	`   �  

  �  

  �  	`   �  	`      B  , ,���  	`���  

����  

����  	`���  	`      B  , ,���+  	`���+  

����  

����  	`���+  	`      B  , ,����  	`����  

����  

����  	`����  	`      B  , ,  �    �  �  5  �  5    �        B  , ,  �    �  �  U  �  U    �        B  , ,  �    �  �  u  �  u    �        B  , ,   �     �  �  �  �  �     �        B  , ,���  ���  �����  �����  ���        B  , ,���+  ���+  �����  �����  ���+        B  , ,����  ����  �����  �����  ����        B  , ,  k  �  k  b  	  b  	  �  k  �      B  , ,  �  �  �  b  5  b  5  �  �  �      B  , ,  �  �  �  b  U  b  U  �  �  �      B  , ,  �  �  �  b  u  b  u  �  �  �      B  , ,   �  �   �  b  �  b  �  �   �  �      B  , ,���  ����  b����  b����  ����  �      B  , ,���+  ����+  b����  b����  ����+  �      B  , ,����  �����  b����  b����  �����  �      B  , ,  k  d  k    	    	  d  k  d      B  , ,  �  d  �    5    5  d  �  d      B  , ,  �  d  �    U    U  d  �  d      B  , ,  �  d  �    u    u  d  �  d      B  , ,   �  d   �    �    �  d   �  d      B  , ,���  d���  ����  ����  d���  d      B  , ,���+  d���+  ����  ����  d���+  d      B  , ,����  d����  ����  ����  d����  d      B  , ,����  ����  �����  �����  ����        B  , ,  k    k  �  	  �  	    k        B  , ,  _���@  _����  	����  	���@  _���@      B  , ,  ���@  ����  �����  ����@  ���@      B  , ,  ����@  �����  a����  a���@  ����@      B  , ,  c���@  c����  ����  ���@  c���@      B  , ,   ���@   ����   �����   ����@   ���@      B  , ,�������@�����������e�������e���@�������@      B  , ,���g���@���g�����������������@���g���@      B  , ,���������������j�������j����������������      B  , ,  k���  k����  	����  	���  k���      B  , ,  ����  �����  5����  5���  ����      B  , ,  ����  �����  U����  U���  ����      B  , ,  ����  �����  u����  u���  ����      B  , ,   ����   �����  �����  ����   ����      B  , ,����������������������������������      B  , ,���+������+����������������������+���      B  , ,�������������������������������������      B  , ,  k���h  k���  	���  	���h  k���h      B  , ,  ����h  ����  5���  5���h  ����h      B  , ,  ����h  ����  U���  U���h  ����h      B  , ,  ����h  ����  u���  u���h  ����h      B  , ,   ����h   ����  ����  ����h   ����h      B  , ,������h��������������������h������h      B  , ,���+���h���+�����������������h���+���h      B  , ,�������h���������������������h�������h      B  , ,���+�������+���f�������f�����������+����      B  , ,���������������f�������f����������������      B  , ,  k  �  k  b  	  b  	  �  k  �      B  , ,  �  �  �  b  5  b  5  �  �  �      B  , ,  �  �  �  b  U  b  U  �  �  �      B  , ,  �  �  �  b  u  b  u  �  �  �      B  , ,   �  �   �  b  �  b  �  �   �  �      B  , ,���  ����  b����  b����  ����  �      B  , ,���+  ����+  b����  b����  ����+  �      B  , ,����  �����  b����  b����  �����  �      B  , ,  k���  k����  	����  	���  k���      B  , ,  ����  �����  5����  5���  ����      B  , ,  ����  �����  U����  U���  ����      B  , ,  ����  �����  u����  u���  ����      B  , ,   ����   �����  �����  ����   ����      B  , ,����������������������������������      B  , ,���+������+����������������������+���      B  , ,�������������������������������������      B  , ,���+   d���+  ����  ����   d���+   d      B  , ,����   d����  ����  ����   d����   d      B  , ,  k����  k���f  	���f  	����  k����      B  , ,  �����  ����f  5���f  5����  �����      B  , ,  �����  ����f  U���f  U����  �����      B  , ,  �����  ����f  u���f  u����  �����      B  , ,   �����   ����f  ����f  �����   �����      B  , ,�������������f�������f���������������      B  , ,  k   d  k    	    	   d  k   d      B  , ,  �   d  �    5    5   d  �   d      B  , ,  �   d  �    U    U   d  �   d      B  , ,  �   d  �    u    u   d  �   d      B  , ,   �   d   �    �    �   d   �   d      B  , ,���   d���  ����  ����   d���   d      B  , ,  ���@  ����  �����  ����@  ���@      B  , ,  ����@  �����  ]����  ]���@  ����@      B  , ,  O���@  O����  �����  ����@  O���@      B  , ,  �  �  �  b  5  b  5  �  �  �      B  , ,  �  �  �  b  U  b  U  �  �  �      B  , ,  �  �  �  b  u  b  u  �  �  �      B  , ,  �  �  �  b  �  b  �  �  �  �      B  , ,    �    b  �  b  �  �    �      B  , ,  
K����  
K���f  
����f  
�����  
K����      B  , ,  ����  �����  o����  o���  ����      B  , ,  ����  �����  5����  5���  ����      B  , ,  ����  �����  U����  U���  ����      B  , ,  ����  �����  u����  u���  ����      B  , ,  ����  �����  �����  ����  ����      B  , ,  ���  ����  �����  ����  ���      B  , ,  +���  +����  �����  ����  +���      B  , ,  
K���  
K����  
�����  
����  
K���      B  , ,  �   d  �    o    o   d  �   d      B  , ,  �   d  �    5    5   d  �   d      B  , ,  �   d  �    U    U   d  �   d      B  , ,  �   d  �    u    u   d  �   d      B  , ,  �   d  �    �    �   d  �   d      B  , ,     d      �    �   d     d      B  , ,  +   d  +    �    �   d  +   d      B  , ,  
K   d  
K    
�    
�   d  
K   d      B  , ,  +���  +����  �����  ����  +���      B  , ,  
K���  
K����  
�����  
����  
K���      B  , ,  +  �  +  b  �  b  �  �  +  �      B  , ,  
K  �  
K  b  
�  b  
�  �  
K  �      B  , ,  �����  ����f  o���f  o����  �����      B  , ,  �����  ����f  5���f  5����  �����      B  , ,  �����  ����f  U���f  U����  �����      B  , ,  �����  ����f  u���f  u����  �����      B  , ,  �����  ����f  ����f  �����  �����      B  , ,  ����  ���f  ����f  �����  ����      B  , ,  +����  +���f  ����f  �����  +����      B  , ,  ����h  ����  o���  o���h  ����h      B  , ,  ����h  ����  5���  5���h  ����h      B  , ,  ����h  ����  U���  U���h  ����h      B  , ,  ����h  ����  u���  u���h  ����h      B  , ,  ����h  ����  ����  ����h  ����h      B  , ,  ���h  ���  ����  ����h  ���h      B  , ,  +���h  +���  ����  ����h  +���h      B  , ,  
K���h  
K���  
����  
����h  
K���h      B  , ,  �����  ����j  o���j  o����  �����      B  , ,  ����@  �����  �����  ����@  ����@      B  , ,  ����  �����  o����  o���  ����      B  , ,  ����  �����  5����  5���  ����      B  , ,  ����  �����  U����  U���  ����      B  , ,  ����  �����  u����  u���  ����      B  , ,  ����  �����  �����  ����  ����      B  , ,  ���  ����  �����  ����  ���      B  , ,  �    �  �  o  �  o    �        B  , ,  �  �  �  b  o  b  o  �  �  �      B  , ,  ����@  �����  Q����  Q���@  ����@      B  , ,  S���@  S����  �����  ����@  S���@      B  , ,  ����@  �����  �����  ����@  ����@      B  , ,  ����@  �����  U����  U���@  ����@      B  , ,  W���@  W����  ����  ���@  W���@      B  , ,  ���@  ����  �����  ����@  ���@      B  , ,  
����@  
�����  Y����  Y���@  
����@      @   ,���=�������=  :  #  :  #�������=����      A   ,������������  �  q  �  q������������      A   ,����  #����  �  q  �  q  #����  #      ]  , ,���t�������t���g  ����g  ��������t����      ]  , ,  H���g  H  _  �  _  ����g  H���g      ]  , ,���t���g���t  _���  _������g���t���g      ]  , ,���t  _���t    �    �  _���t  _     �     0�     0 mimcap_1    F   ,              >�  @o  >�  @o                  G   ,  �  �  �  ;�  ;�  ;�  ;�  �  �  �      G   ,  >{   <  >{  >D  @[  >D  @[   <  >{   <      F  , ,  !4  �  !4  L  !�  L  !�  �  !4  �      F  , ,  !4  �  !4  L  !�  L  !�  �  !4  �      F  , ,  !4    !4  �  !�  �  !�    !4        F  , ,  !4    !4  �  !�  �  !�    !4        F  , ,  !4  �  !4  l  !�  l  !�  �  !4  �      F  , ,  !4  �  !4  l  !�  l  !�  �  !4  �      F  , ,  !4  4  !4  �  !�  �  !�  4  !4  4      F  , ,  !4  4  !4  �  !�  �  !�  4  !4  4      F  , ,  !4  	�  !4  
�  !�  
�  !�  	�  !4  	�      F  , ,  !4  	�  !4  
�  !�  
�  !�  	�  !4  	�      F  , ,  !4  T  !4    !�    !�  T  !4  T      F  , ,  !4  T  !4    !�    !�  T  !4  T      F  , ,  !4  �  !4  �  !�  �  !�  �  !4  �      F  , ,  !4  �  !4  �  !�  �  !�  �  !4  �      F  , ,  !4  t  !4  <  !�  <  !�  t  !4  t      F  , ,  !4  t  !4  <  !�  <  !�  t  !4  t      F  , ,  !4    !4  �  !�  �  !�    !4        F  , ,  !4    !4  �  !�  �  !�    !4        F  , ,  !4  �  !4  \  !�  \  !�  �  !4  �      F  , ,  !4  �  !4  \  !�  \  !�  �  !4  �      F  , ,  !4  $  !4  �  !�  �  !�  $  !4  $      F  , ,  !4  $  !4  �  !�  �  !�  $  !4  $      F  , ,  !4  �  !4  |  !�  |  !�  �  !4  �      F  , ,  !4  �  !4  |  !�  |  !�  �  !4  �      F  , ,  !4  D  !4    !�    !�  D  !4  D      F  , ,  !4  D  !4    !�    !�  D  !4  D      F  , ,  !4  �  !4  �  !�  �  !�  �  !4  �      F  , ,  !4  �  !4  �  !�  �  !�  �  !4  �      F  , ,  !4  d  !4  ,  !�  ,  !�  d  !4  d      F  , ,  !4  d  !4  ,  !�  ,  !�  d  !4  d      F  , ,  !4  �  !4  �  !�  �  !�  �  !4  �      F  , ,  !4  �  !4  �  !�  �  !�  �  !4  �      F  , ,  !4  �  !4  L  !�  L  !�  �  !4  �      F  , ,  !4  �  !4  L  !�  L  !�  �  !4  �      F  , ,  !4    !4  �  !�  �  !�    !4        F  , ,  !4    !4  �  !�  �  !�    !4        F  , ,  !4  �  !4   l  !�   l  !�  �  !4  �      F  , ,  !4  �  !4   l  !�   l  !�  �  !4  �      F  , ,  !4  !4  !4  !�  !�  !�  !�  !4  !4  !4      F  , ,  !4  !4  !4  !�  !�  !�  !�  !4  !4  !4      F  , ,  !4  "�  !4  #�  !�  #�  !�  "�  !4  "�      F  , ,  !4  "�  !4  #�  !�  #�  !�  "�  !4  "�      F  , ,  !4  $T  !4  %  !�  %  !�  $T  !4  $T      F  , ,  !4  $T  !4  %  !�  %  !�  $T  !4  $T      F  , ,  !4  %�  !4  &�  !�  &�  !�  %�  !4  %�      F  , ,  !4  %�  !4  &�  !�  &�  !�  %�  !4  %�      F  , ,  !4  't  !4  (<  !�  (<  !�  't  !4  't      F  , ,  !4  't  !4  (<  !�  (<  !�  't  !4  't      F  , ,  !4  )  !4  )�  !�  )�  !�  )  !4  )      F  , ,  !4  )  !4  )�  !�  )�  !�  )  !4  )      F  , ,  !4  *�  !4  +\  !�  +\  !�  *�  !4  *�      F  , ,  !4  *�  !4  +\  !�  +\  !�  *�  !4  *�      F  , ,  !4  ,$  !4  ,�  !�  ,�  !�  ,$  !4  ,$      F  , ,  !4  ,$  !4  ,�  !�  ,�  !�  ,$  !4  ,$      F  , ,  !4  -�  !4  .|  !�  .|  !�  -�  !4  -�      F  , ,  !4  -�  !4  .|  !�  .|  !�  -�  !4  -�      F  , ,  !4  /D  !4  0  !�  0  !�  /D  !4  /D      F  , ,  !4  /D  !4  0  !�  0  !�  /D  !4  /D      F  , ,  !4  0�  !4  1�  !�  1�  !�  0�  !4  0�      F  , ,  !4  0�  !4  1�  !�  1�  !�  0�  !4  0�      F  , ,  !4  2d  !4  3,  !�  3,  !�  2d  !4  2d      F  , ,  !4  2d  !4  3,  !�  3,  !�  2d  !4  2d      F  , ,  !4  3�  !4  4�  !�  4�  !�  3�  !4  3�      F  , ,  !4  3�  !4  4�  !�  4�  !�  3�  !4  3�      F  , ,  !4  5�  !4  6L  !�  6L  !�  5�  !4  5�      F  , ,  !4  5�  !4  6L  !�  6L  !�  5�  !4  5�      F  , ,  !4  7  !4  7�  !�  7�  !�  7  !4  7      F  , ,  !4  7  !4  7�  !�  7�  !�  7  !4  7      F  , ,  !4  8�  !4  9l  !�  9l  !�  8�  !4  8�      F  , ,  !4  8�  !4  9l  !�  9l  !�  8�  !4  8�      F  , ,  !4  :4  !4  :�  !�  :�  !�  :4  !4  :4      F  , ,  !4  :4  !4  :�  !�  :�  !�  :4  !4  :4      F  , ,  ?  �  ?  �  ?�  �  ?�  �  ?  �      F  , ,  ?  �  ?  �  ?�  �  ?�  �  ?  �      F  , ,  "�  -�  "�  .|  #�  .|  #�  -�  "�  -�      F  , ,  "�  -�  "�  .|  #�  .|  #�  -�  "�  -�      F  , ,  $T  -�  $T  .|  %  .|  %  -�  $T  -�      F  , ,  $T  -�  $T  .|  %  .|  %  -�  $T  -�      F  , ,  %�  -�  %�  .|  &�  .|  &�  -�  %�  -�      F  , ,  %�  -�  %�  .|  &�  .|  &�  -�  %�  -�      F  , ,  't  -�  't  .|  (<  .|  (<  -�  't  -�      F  , ,  't  -�  't  .|  (<  .|  (<  -�  't  -�      F  , ,  )  -�  )  .|  )�  .|  )�  -�  )  -�      F  , ,  )  -�  )  .|  )�  .|  )�  -�  )  -�      F  , ,  *�  -�  *�  .|  +\  .|  +\  -�  *�  -�      F  , ,  *�  -�  *�  .|  +\  .|  +\  -�  *�  -�      F  , ,  ,$  -�  ,$  .|  ,�  .|  ,�  -�  ,$  -�      F  , ,  ,$  -�  ,$  .|  ,�  .|  ,�  -�  ,$  -�      F  , ,  -�  -�  -�  .|  .|  .|  .|  -�  -�  -�      F  , ,  -�  -�  -�  .|  .|  .|  .|  -�  -�  -�      F  , ,  /D  -�  /D  .|  0  .|  0  -�  /D  -�      F  , ,  /D  -�  /D  .|  0  .|  0  -�  /D  -�      F  , ,  0�  -�  0�  .|  1�  .|  1�  -�  0�  -�      F  , ,  0�  -�  0�  .|  1�  .|  1�  -�  0�  -�      F  , ,  2d  -�  2d  .|  3,  .|  3,  -�  2d  -�      F  , ,  2d  -�  2d  .|  3,  .|  3,  -�  2d  -�      F  , ,  3�  -�  3�  .|  4�  .|  4�  -�  3�  -�      F  , ,  3�  -�  3�  .|  4�  .|  4�  -�  3�  -�      F  , ,  5�  -�  5�  .|  6L  .|  6L  -�  5�  -�      F  , ,  5�  -�  5�  .|  6L  .|  6L  -�  5�  -�      F  , ,  7  -�  7  .|  7�  .|  7�  -�  7  -�      F  , ,  7  -�  7  .|  7�  .|  7�  -�  7  -�      F  , ,  8�  -�  8�  .|  9l  .|  9l  -�  8�  -�      F  , ,  8�  -�  8�  .|  9l  .|  9l  -�  8�  -�      F  , ,  :4  -�  :4  .|  :�  .|  :�  -�  :4  -�      F  , ,  :4  -�  :4  .|  :�  .|  :�  -�  :4  -�      F  , ,  0�  5�  0�  6L  1�  6L  1�  5�  0�  5�      F  , ,  0�  5�  0�  6L  1�  6L  1�  5�  0�  5�      F  , ,  2d  5�  2d  6L  3,  6L  3,  5�  2d  5�      F  , ,  2d  5�  2d  6L  3,  6L  3,  5�  2d  5�      F  , ,  3�  5�  3�  6L  4�  6L  4�  5�  3�  5�      F  , ,  3�  5�  3�  6L  4�  6L  4�  5�  3�  5�      F  , ,  5�  5�  5�  6L  6L  6L  6L  5�  5�  5�      F  , ,  5�  5�  5�  6L  6L  6L  6L  5�  5�  5�      F  , ,  7  5�  7  6L  7�  6L  7�  5�  7  5�      F  , ,  7  5�  7  6L  7�  6L  7�  5�  7  5�      F  , ,  8�  5�  8�  6L  9l  6L  9l  5�  8�  5�      F  , ,  8�  5�  8�  6L  9l  6L  9l  5�  8�  5�      F  , ,  :4  5�  :4  6L  :�  6L  :�  5�  :4  5�      F  , ,  :4  5�  :4  6L  :�  6L  :�  5�  :4  5�      F  , ,  8�  7  8�  7�  9l  7�  9l  7  8�  7      F  , ,  8�  7  8�  7�  9l  7�  9l  7  8�  7      F  , ,  :4  7  :4  7�  :�  7�  :�  7  :4  7      F  , ,  :4  7  :4  7�  :�  7�  :�  7  :4  7      F  , ,  8�  8�  8�  9l  9l  9l  9l  8�  8�  8�      F  , ,  8�  8�  8�  9l  9l  9l  9l  8�  8�  8�      F  , ,  :4  8�  :4  9l  :�  9l  :�  8�  :4  8�      F  , ,  :4  8�  :4  9l  :�  9l  :�  8�  :4  8�      F  , ,  8�  :4  8�  :�  9l  :�  9l  :4  8�  :4      F  , ,  8�  :4  8�  :�  9l  :�  9l  :4  8�  :4      F  , ,  :4  :4  :4  :�  :�  :�  :�  :4  :4  :4      F  , ,  :4  :4  :4  :�  :�  :�  :�  :4  :4  :4      F  , ,  ?  6L  ?  7  ?�  7  ?�  6L  ?  6L      F  , ,  ?  6L  ?  7  ?�  7  ?�  6L  ?  6L      F  , ,  ?  7�  ?  8�  ?�  8�  ?�  7�  ?  7�      F  , ,  ?  7�  ?  8�  ?�  8�  ?�  7�  ?  7�      F  , ,  ?  9l  ?  :4  ?�  :4  ?�  9l  ?  9l      F  , ,  ?  9l  ?  :4  ?�  :4  ?�  9l  ?  9l      F  , ,  ?  :�  ?  ;�  ?�  ;�  ?�  :�  ?  :�      F  , ,  ?  :�  ?  ;�  ?�  ;�  ?�  :�  ?  :�      F  , ,  ?  <�  ?  =T  ?�  =T  ?�  <�  ?  <�      F  , ,  ?  <�  ?  =T  ?�  =T  ?�  <�  ?  <�      F  , ,  7  8�  7  9l  7�  9l  7�  8�  7  8�      F  , ,  7  8�  7  9l  7�  9l  7�  8�  7  8�      F  , ,  3�  7  3�  7�  4�  7�  4�  7  3�  7      F  , ,  3�  7  3�  7�  4�  7�  4�  7  3�  7      F  , ,  5�  7  5�  7�  6L  7�  6L  7  5�  7      F  , ,  5�  7  5�  7�  6L  7�  6L  7  5�  7      F  , ,  0�  :4  0�  :�  1�  :�  1�  :4  0�  :4      F  , ,  0�  :4  0�  :�  1�  :�  1�  :4  0�  :4      F  , ,  2d  :4  2d  :�  3,  :�  3,  :4  2d  :4      F  , ,  2d  :4  2d  :�  3,  :�  3,  :4  2d  :4      F  , ,  3�  :4  3�  :�  4�  :�  4�  :4  3�  :4      F  , ,  3�  :4  3�  :�  4�  :�  4�  :4  3�  :4      F  , ,  5�  :4  5�  :�  6L  :�  6L  :4  5�  :4      F  , ,  5�  :4  5�  :�  6L  :�  6L  :4  5�  :4      F  , ,  7  :4  7  :�  7�  :�  7�  :4  7  :4      F  , ,  7  :4  7  :�  7�  :�  7�  :4  7  :4      F  , ,  7  7  7  7�  7�  7�  7�  7  7  7      F  , ,  7  7  7  7�  7�  7�  7�  7  7  7      F  , ,  0�  7  0�  7�  1�  7�  1�  7  0�  7      F  , ,  0�  7  0�  7�  1�  7�  1�  7  0�  7      F  , ,  2d  7  2d  7�  3,  7�  3,  7  2d  7      F  , ,  2d  7  2d  7�  3,  7�  3,  7  2d  7      F  , ,  0�  8�  0�  9l  1�  9l  1�  8�  0�  8�      F  , ,  0�  8�  0�  9l  1�  9l  1�  8�  0�  8�      F  , ,  2d  8�  2d  9l  3,  9l  3,  8�  2d  8�      F  , ,  2d  8�  2d  9l  3,  9l  3,  8�  2d  8�      F  , ,  3�  8�  3�  9l  4�  9l  4�  8�  3�  8�      F  , ,  3�  8�  3�  9l  4�  9l  4�  8�  3�  8�      F  , ,  5�  8�  5�  9l  6L  9l  6L  8�  5�  8�      F  , ,  5�  8�  5�  9l  6L  9l  6L  8�  5�  8�      F  , ,  5�  2d  5�  3,  6L  3,  6L  2d  5�  2d      F  , ,  5�  2d  5�  3,  6L  3,  6L  2d  5�  2d      F  , ,  7  2d  7  3,  7�  3,  7�  2d  7  2d      F  , ,  7  2d  7  3,  7�  3,  7�  2d  7  2d      F  , ,  0�  3�  0�  4�  1�  4�  1�  3�  0�  3�      F  , ,  0�  3�  0�  4�  1�  4�  1�  3�  0�  3�      F  , ,  2d  3�  2d  4�  3,  4�  3,  3�  2d  3�      F  , ,  2d  3�  2d  4�  3,  4�  3,  3�  2d  3�      F  , ,  3�  3�  3�  4�  4�  4�  4�  3�  3�  3�      F  , ,  3�  3�  3�  4�  4�  4�  4�  3�  3�  3�      F  , ,  5�  3�  5�  4�  6L  4�  6L  3�  5�  3�      F  , ,  5�  3�  5�  4�  6L  4�  6L  3�  5�  3�      F  , ,  7  3�  7  4�  7�  4�  7�  3�  7  3�      F  , ,  7  3�  7  4�  7�  4�  7�  3�  7  3�      F  , ,  0�  /D  0�  0  1�  0  1�  /D  0�  /D      F  , ,  0�  /D  0�  0  1�  0  1�  /D  0�  /D      F  , ,  2d  /D  2d  0  3,  0  3,  /D  2d  /D      F  , ,  2d  /D  2d  0  3,  0  3,  /D  2d  /D      F  , ,  3�  /D  3�  0  4�  0  4�  /D  3�  /D      F  , ,  3�  /D  3�  0  4�  0  4�  /D  3�  /D      F  , ,  5�  /D  5�  0  6L  0  6L  /D  5�  /D      F  , ,  5�  /D  5�  0  6L  0  6L  /D  5�  /D      F  , ,  7  /D  7  0  7�  0  7�  /D  7  /D      F  , ,  7  /D  7  0  7�  0  7�  /D  7  /D      F  , ,  0�  0�  0�  1�  1�  1�  1�  0�  0�  0�      F  , ,  0�  0�  0�  1�  1�  1�  1�  0�  0�  0�      F  , ,  2d  0�  2d  1�  3,  1�  3,  0�  2d  0�      F  , ,  2d  0�  2d  1�  3,  1�  3,  0�  2d  0�      F  , ,  3�  0�  3�  1�  4�  1�  4�  0�  3�  0�      F  , ,  3�  0�  3�  1�  4�  1�  4�  0�  3�  0�      F  , ,  5�  0�  5�  1�  6L  1�  6L  0�  5�  0�      F  , ,  5�  0�  5�  1�  6L  1�  6L  0�  5�  0�      F  , ,  7  0�  7  1�  7�  1�  7�  0�  7  0�      F  , ,  7  0�  7  1�  7�  1�  7�  0�  7  0�      F  , ,  0�  2d  0�  3,  1�  3,  1�  2d  0�  2d      F  , ,  0�  2d  0�  3,  1�  3,  1�  2d  0�  2d      F  , ,  2d  2d  2d  3,  3,  3,  3,  2d  2d  2d      F  , ,  2d  2d  2d  3,  3,  3,  3,  2d  2d  2d      F  , ,  3�  2d  3�  3,  4�  3,  4�  2d  3�  2d      F  , ,  3�  2d  3�  3,  4�  3,  4�  2d  3�  2d      F  , ,  8�  /D  8�  0  9l  0  9l  /D  8�  /D      F  , ,  8�  /D  8�  0  9l  0  9l  /D  8�  /D      F  , ,  8�  0�  8�  1�  9l  1�  9l  0�  8�  0�      F  , ,  8�  0�  8�  1�  9l  1�  9l  0�  8�  0�      F  , ,  :4  0�  :4  1�  :�  1�  :�  0�  :4  0�      F  , ,  :4  0�  :4  1�  :�  1�  :�  0�  :4  0�      F  , ,  ?  .|  ?  /D  ?�  /D  ?�  .|  ?  .|      F  , ,  ?  .|  ?  /D  ?�  /D  ?�  .|  ?  .|      F  , ,  ?  0  ?  0�  ?�  0�  ?�  0  ?  0      F  , ,  ?  0  ?  0�  ?�  0�  ?�  0  ?  0      F  , ,  ?  1�  ?  2d  ?�  2d  ?�  1�  ?  1�      F  , ,  ?  1�  ?  2d  ?�  2d  ?�  1�  ?  1�      F  , ,  ?  3,  ?  3�  ?�  3�  ?�  3,  ?  3,      F  , ,  ?  3,  ?  3�  ?�  3�  ?�  3,  ?  3,      F  , ,  ?  4�  ?  5�  ?�  5�  ?�  4�  ?  4�      F  , ,  ?  4�  ?  5�  ?�  5�  ?�  4�  ?  4�      F  , ,  :4  /D  :4  0  :�  0  :�  /D  :4  /D      F  , ,  :4  /D  :4  0  :�  0  :�  /D  :4  /D      F  , ,  8�  2d  8�  3,  9l  3,  9l  2d  8�  2d      F  , ,  8�  2d  8�  3,  9l  3,  9l  2d  8�  2d      F  , ,  8�  3�  8�  4�  9l  4�  9l  3�  8�  3�      F  , ,  8�  3�  8�  4�  9l  4�  9l  3�  8�  3�      F  , ,  :4  3�  :4  4�  :�  4�  :�  3�  :4  3�      F  , ,  :4  3�  :4  4�  :�  4�  :�  3�  :4  3�      F  , ,  :4  2d  :4  3,  :�  3,  :�  2d  :4  2d      F  , ,  :4  2d  :4  3,  :�  3,  :�  2d  :4  2d      F  , ,  %�  5�  %�  6L  &�  6L  &�  5�  %�  5�      F  , ,  %�  5�  %�  6L  &�  6L  &�  5�  %�  5�      F  , ,  't  5�  't  6L  (<  6L  (<  5�  't  5�      F  , ,  't  5�  't  6L  (<  6L  (<  5�  't  5�      F  , ,  )  5�  )  6L  )�  6L  )�  5�  )  5�      F  , ,  )  5�  )  6L  )�  6L  )�  5�  )  5�      F  , ,  *�  5�  *�  6L  +\  6L  +\  5�  *�  5�      F  , ,  *�  5�  *�  6L  +\  6L  +\  5�  *�  5�      F  , ,  ,$  5�  ,$  6L  ,�  6L  ,�  5�  ,$  5�      F  , ,  ,$  5�  ,$  6L  ,�  6L  ,�  5�  ,$  5�      F  , ,  -�  5�  -�  6L  .|  6L  .|  5�  -�  5�      F  , ,  -�  5�  -�  6L  .|  6L  .|  5�  -�  5�      F  , ,  /D  5�  /D  6L  0  6L  0  5�  /D  5�      F  , ,  /D  5�  /D  6L  0  6L  0  5�  /D  5�      F  , ,  )  /D  )  0  )�  0  )�  /D  )  /D      F  , ,  )  /D  )  0  )�  0  )�  /D  )  /D      F  , ,  )  7  )  7�  )�  7�  )�  7  )  7      F  , ,  )  7  )  7�  )�  7�  )�  7  )  7      F  , ,  )  2d  )  3,  )�  3,  )�  2d  )  2d      F  , ,  )  2d  )  3,  )�  3,  )�  2d  )  2d      F  , ,  )  8�  )  9l  )�  9l  )�  8�  )  8�      F  , ,  )  8�  )  9l  )�  9l  )�  8�  )  8�      F  , ,  )  0�  )  1�  )�  1�  )�  0�  )  0�      F  , ,  )  0�  )  1�  )�  1�  )�  0�  )  0�      F  , ,  )  :4  )  :�  )�  :�  )�  :4  )  :4      F  , ,  )  :4  )  :�  )�  :�  )�  :4  )  :4      F  , ,  )  3�  )  4�  )�  4�  )�  3�  )  3�      F  , ,  )  3�  )  4�  )�  4�  )�  3�  )  3�      F  , ,  "�  5�  "�  6L  #�  6L  #�  5�  "�  5�      F  , ,  "�  5�  "�  6L  #�  6L  #�  5�  "�  5�      F  , ,  $T  5�  $T  6L  %  6L  %  5�  $T  5�      F  , ,  $T  5�  $T  6L  %  6L  %  5�  $T  5�      F  , ,  ,$  8�  ,$  9l  ,�  9l  ,�  8�  ,$  8�      F  , ,  ,$  8�  ,$  9l  ,�  9l  ,�  8�  ,$  8�      F  , ,  -�  8�  -�  9l  .|  9l  .|  8�  -�  8�      F  , ,  -�  8�  -�  9l  .|  9l  .|  8�  -�  8�      F  , ,  /D  8�  /D  9l  0  9l  0  8�  /D  8�      F  , ,  /D  8�  /D  9l  0  9l  0  8�  /D  8�      F  , ,  -�  7  -�  7�  .|  7�  .|  7  -�  7      F  , ,  -�  7  -�  7�  .|  7�  .|  7  -�  7      F  , ,  /D  7  /D  7�  0  7�  0  7  /D  7      F  , ,  /D  7  /D  7�  0  7�  0  7  /D  7      F  , ,  *�  :4  *�  :�  +\  :�  +\  :4  *�  :4      F  , ,  *�  :4  *�  :�  +\  :�  +\  :4  *�  :4      F  , ,  ,$  :4  ,$  :�  ,�  :�  ,�  :4  ,$  :4      F  , ,  ,$  :4  ,$  :�  ,�  :�  ,�  :4  ,$  :4      F  , ,  -�  :4  -�  :�  .|  :�  .|  :4  -�  :4      F  , ,  -�  :4  -�  :�  .|  :�  .|  :4  -�  :4      F  , ,  /D  :4  /D  :�  0  :�  0  :4  /D  :4      F  , ,  /D  :4  /D  :�  0  :�  0  :4  /D  :4      F  , ,  *�  7  *�  7�  +\  7�  +\  7  *�  7      F  , ,  *�  7  *�  7�  +\  7�  +\  7  *�  7      F  , ,  ,$  7  ,$  7�  ,�  7�  ,�  7  ,$  7      F  , ,  ,$  7  ,$  7�  ,�  7�  ,�  7  ,$  7      F  , ,  *�  8�  *�  9l  +\  9l  +\  8�  *�  8�      F  , ,  *�  8�  *�  9l  +\  9l  +\  8�  *�  8�      F  , ,  "�  :4  "�  :�  #�  :�  #�  :4  "�  :4      F  , ,  "�  :4  "�  :�  #�  :�  #�  :4  "�  :4      F  , ,  $T  :4  $T  :�  %  :�  %  :4  $T  :4      F  , ,  $T  :4  $T  :�  %  :�  %  :4  $T  :4      F  , ,  %�  :4  %�  :�  &�  :�  &�  :4  %�  :4      F  , ,  %�  :4  %�  :�  &�  :�  &�  :4  %�  :4      F  , ,  't  :4  't  :�  (<  :�  (<  :4  't  :4      F  , ,  't  :4  't  :�  (<  :�  (<  :4  't  :4      F  , ,  %�  8�  %�  9l  &�  9l  &�  8�  %�  8�      F  , ,  %�  8�  %�  9l  &�  9l  &�  8�  %�  8�      F  , ,  't  8�  't  9l  (<  9l  (<  8�  't  8�      F  , ,  't  8�  't  9l  (<  9l  (<  8�  't  8�      F  , ,  %�  7  %�  7�  &�  7�  &�  7  %�  7      F  , ,  %�  7  %�  7�  &�  7�  &�  7  %�  7      F  , ,  't  7  't  7�  (<  7�  (<  7  't  7      F  , ,  't  7  't  7�  (<  7�  (<  7  't  7      F  , ,  "�  7  "�  7�  #�  7�  #�  7  "�  7      F  , ,  "�  7  "�  7�  #�  7�  #�  7  "�  7      F  , ,  $T  7  $T  7�  %  7�  %  7  $T  7      F  , ,  $T  7  $T  7�  %  7�  %  7  $T  7      F  , ,  "�  8�  "�  9l  #�  9l  #�  8�  "�  8�      F  , ,  "�  8�  "�  9l  #�  9l  #�  8�  "�  8�      F  , ,  $T  8�  $T  9l  %  9l  %  8�  $T  8�      F  , ,  $T  8�  $T  9l  %  9l  %  8�  $T  8�      F  , ,  't  /D  't  0  (<  0  (<  /D  't  /D      F  , ,  't  /D  't  0  (<  0  (<  /D  't  /D      F  , ,  $T  /D  $T  0  %  0  %  /D  $T  /D      F  , ,  $T  /D  $T  0  %  0  %  /D  $T  /D      F  , ,  't  2d  't  3,  (<  3,  (<  2d  't  2d      F  , ,  't  2d  't  3,  (<  3,  (<  2d  't  2d      F  , ,  "�  2d  "�  3,  #�  3,  #�  2d  "�  2d      F  , ,  "�  2d  "�  3,  #�  3,  #�  2d  "�  2d      F  , ,  $T  2d  $T  3,  %  3,  %  2d  $T  2d      F  , ,  $T  2d  $T  3,  %  3,  %  2d  $T  2d      F  , ,  %�  2d  %�  3,  &�  3,  &�  2d  %�  2d      F  , ,  %�  2d  %�  3,  &�  3,  &�  2d  %�  2d      F  , ,  "�  0�  "�  1�  #�  1�  #�  0�  "�  0�      F  , ,  "�  0�  "�  1�  #�  1�  #�  0�  "�  0�      F  , ,  $T  0�  $T  1�  %  1�  %  0�  $T  0�      F  , ,  $T  0�  $T  1�  %  1�  %  0�  $T  0�      F  , ,  %�  0�  %�  1�  &�  1�  &�  0�  %�  0�      F  , ,  %�  0�  %�  1�  &�  1�  &�  0�  %�  0�      F  , ,  $T  3�  $T  4�  %  4�  %  3�  $T  3�      F  , ,  $T  3�  $T  4�  %  4�  %  3�  $T  3�      F  , ,  %�  3�  %�  4�  &�  4�  &�  3�  %�  3�      F  , ,  %�  3�  %�  4�  &�  4�  &�  3�  %�  3�      F  , ,  't  3�  't  4�  (<  4�  (<  3�  't  3�      F  , ,  't  3�  't  4�  (<  4�  (<  3�  't  3�      F  , ,  't  0�  't  1�  (<  1�  (<  0�  't  0�      F  , ,  't  0�  't  1�  (<  1�  (<  0�  't  0�      F  , ,  "�  /D  "�  0  #�  0  #�  /D  "�  /D      F  , ,  "�  /D  "�  0  #�  0  #�  /D  "�  /D      F  , ,  %�  /D  %�  0  &�  0  &�  /D  %�  /D      F  , ,  %�  /D  %�  0  &�  0  &�  /D  %�  /D      F  , ,  "�  3�  "�  4�  #�  4�  #�  3�  "�  3�      F  , ,  "�  3�  "�  4�  #�  4�  #�  3�  "�  3�      F  , ,  /D  2d  /D  3,  0  3,  0  2d  /D  2d      F  , ,  /D  2d  /D  3,  0  3,  0  2d  /D  2d      F  , ,  ,$  /D  ,$  0  ,�  0  ,�  /D  ,$  /D      F  , ,  ,$  /D  ,$  0  ,�  0  ,�  /D  ,$  /D      F  , ,  *�  /D  *�  0  +\  0  +\  /D  *�  /D      F  , ,  *�  /D  *�  0  +\  0  +\  /D  *�  /D      F  , ,  *�  3�  *�  4�  +\  4�  +\  3�  *�  3�      F  , ,  *�  3�  *�  4�  +\  4�  +\  3�  *�  3�      F  , ,  ,$  3�  ,$  4�  ,�  4�  ,�  3�  ,$  3�      F  , ,  ,$  3�  ,$  4�  ,�  4�  ,�  3�  ,$  3�      F  , ,  -�  3�  -�  4�  .|  4�  .|  3�  -�  3�      F  , ,  -�  3�  -�  4�  .|  4�  .|  3�  -�  3�      F  , ,  /D  3�  /D  4�  0  4�  0  3�  /D  3�      F  , ,  /D  3�  /D  4�  0  4�  0  3�  /D  3�      F  , ,  *�  0�  *�  1�  +\  1�  +\  0�  *�  0�      F  , ,  *�  0�  *�  1�  +\  1�  +\  0�  *�  0�      F  , ,  ,$  0�  ,$  1�  ,�  1�  ,�  0�  ,$  0�      F  , ,  ,$  0�  ,$  1�  ,�  1�  ,�  0�  ,$  0�      F  , ,  -�  0�  -�  1�  .|  1�  .|  0�  -�  0�      F  , ,  -�  0�  -�  1�  .|  1�  .|  0�  -�  0�      F  , ,  /D  0�  /D  1�  0  1�  0  0�  /D  0�      F  , ,  /D  0�  /D  1�  0  1�  0  0�  /D  0�      F  , ,  -�  /D  -�  0  .|  0  .|  /D  -�  /D      F  , ,  -�  /D  -�  0  .|  0  .|  /D  -�  /D      F  , ,  /D  /D  /D  0  0  0  0  /D  /D  /D      F  , ,  /D  /D  /D  0  0  0  0  /D  /D  /D      F  , ,  *�  2d  *�  3,  +\  3,  +\  2d  *�  2d      F  , ,  *�  2d  *�  3,  +\  3,  +\  2d  *�  2d      F  , ,  ,$  2d  ,$  3,  ,�  3,  ,�  2d  ,$  2d      F  , ,  ,$  2d  ,$  3,  ,�  3,  ,�  2d  ,$  2d      F  , ,  -�  2d  -�  3,  .|  3,  .|  2d  -�  2d      F  , ,  -�  2d  -�  3,  .|  3,  .|  2d  -�  2d      F  , ,  )  !4  )  !�  )�  !�  )�  !4  )  !4      F  , ,  )  !4  )  !�  )�  !�  )�  !4  )  !4      F  , ,  )  "�  )  #�  )�  #�  )�  "�  )  "�      F  , ,  )  "�  )  #�  )�  #�  )�  "�  )  "�      F  , ,  )  $T  )  %  )�  %  )�  $T  )  $T      F  , ,  )  $T  )  %  )�  %  )�  $T  )  $T      F  , ,  )  %�  )  &�  )�  &�  )�  %�  )  %�      F  , ,  )  %�  )  &�  )�  &�  )�  %�  )  %�      F  , ,  )  �  )   l  )�   l  )�  �  )  �      F  , ,  )  �  )   l  )�   l  )�  �  )  �      F  , ,  )  't  )  (<  )�  (<  )�  't  )  't      F  , ,  )  't  )  (<  )�  (<  )�  't  )  't      F  , ,  )  )  )  )�  )�  )�  )�  )  )  )      F  , ,  )  )  )  )�  )�  )�  )�  )  )  )      F  , ,  )  *�  )  +\  )�  +\  )�  *�  )  *�      F  , ,  )  *�  )  +\  )�  +\  )�  *�  )  *�      F  , ,  )  ,$  )  ,�  )�  ,�  )�  ,$  )  ,$      F  , ,  )  ,$  )  ,�  )�  ,�  )�  ,$  )  ,$      F  , ,  *�  't  *�  (<  +\  (<  +\  't  *�  't      F  , ,  *�  't  *�  (<  +\  (<  +\  't  *�  't      F  , ,  ,$  't  ,$  (<  ,�  (<  ,�  't  ,$  't      F  , ,  ,$  't  ,$  (<  ,�  (<  ,�  't  ,$  't      F  , ,  -�  't  -�  (<  .|  (<  .|  't  -�  't      F  , ,  -�  't  -�  (<  .|  (<  .|  't  -�  't      F  , ,  /D  't  /D  (<  0  (<  0  't  /D  't      F  , ,  /D  't  /D  (<  0  (<  0  't  /D  't      F  , ,  ,$  ,$  ,$  ,�  ,�  ,�  ,�  ,$  ,$  ,$      F  , ,  ,$  ,$  ,$  ,�  ,�  ,�  ,�  ,$  ,$  ,$      F  , ,  *�  )  *�  )�  +\  )�  +\  )  *�  )      F  , ,  *�  )  *�  )�  +\  )�  +\  )  *�  )      F  , ,  ,$  )  ,$  )�  ,�  )�  ,�  )  ,$  )      F  , ,  ,$  )  ,$  )�  ,�  )�  ,�  )  ,$  )      F  , ,  -�  )  -�  )�  .|  )�  .|  )  -�  )      F  , ,  -�  )  -�  )�  .|  )�  .|  )  -�  )      F  , ,  /D  )  /D  )�  0  )�  0  )  /D  )      F  , ,  /D  )  /D  )�  0  )�  0  )  /D  )      F  , ,  -�  ,$  -�  ,�  .|  ,�  .|  ,$  -�  ,$      F  , ,  -�  ,$  -�  ,�  .|  ,�  .|  ,$  -�  ,$      F  , ,  *�  *�  *�  +\  +\  +\  +\  *�  *�  *�      F  , ,  *�  *�  *�  +\  +\  +\  +\  *�  *�  *�      F  , ,  ,$  *�  ,$  +\  ,�  +\  ,�  *�  ,$  *�      F  , ,  ,$  *�  ,$  +\  ,�  +\  ,�  *�  ,$  *�      F  , ,  -�  *�  -�  +\  .|  +\  .|  *�  -�  *�      F  , ,  -�  *�  -�  +\  .|  +\  .|  *�  -�  *�      F  , ,  /D  *�  /D  +\  0  +\  0  *�  /D  *�      F  , ,  /D  *�  /D  +\  0  +\  0  *�  /D  *�      F  , ,  /D  ,$  /D  ,�  0  ,�  0  ,$  /D  ,$      F  , ,  /D  ,$  /D  ,�  0  ,�  0  ,$  /D  ,$      F  , ,  *�  ,$  *�  ,�  +\  ,�  +\  ,$  *�  ,$      F  , ,  *�  ,$  *�  ,�  +\  ,�  +\  ,$  *�  ,$      F  , ,  "�  )  "�  )�  #�  )�  #�  )  "�  )      F  , ,  "�  )  "�  )�  #�  )�  #�  )  "�  )      F  , ,  "�  *�  "�  +\  #�  +\  #�  *�  "�  *�      F  , ,  "�  *�  "�  +\  #�  +\  #�  *�  "�  *�      F  , ,  $T  *�  $T  +\  %  +\  %  *�  $T  *�      F  , ,  $T  *�  $T  +\  %  +\  %  *�  $T  *�      F  , ,  %�  *�  %�  +\  &�  +\  &�  *�  %�  *�      F  , ,  %�  *�  %�  +\  &�  +\  &�  *�  %�  *�      F  , ,  't  *�  't  +\  (<  +\  (<  *�  't  *�      F  , ,  't  *�  't  +\  (<  +\  (<  *�  't  *�      F  , ,  $T  )  $T  )�  %  )�  %  )  $T  )      F  , ,  $T  )  $T  )�  %  )�  %  )  $T  )      F  , ,  %�  )  %�  )�  &�  )�  &�  )  %�  )      F  , ,  %�  )  %�  )�  &�  )�  &�  )  %�  )      F  , ,  't  )  't  )�  (<  )�  (<  )  't  )      F  , ,  't  )  't  )�  (<  )�  (<  )  't  )      F  , ,  $T  't  $T  (<  %  (<  %  't  $T  't      F  , ,  $T  't  $T  (<  %  (<  %  't  $T  't      F  , ,  %�  't  %�  (<  &�  (<  &�  't  %�  't      F  , ,  %�  't  %�  (<  &�  (<  &�  't  %�  't      F  , ,  "�  ,$  "�  ,�  #�  ,�  #�  ,$  "�  ,$      F  , ,  "�  ,$  "�  ,�  #�  ,�  #�  ,$  "�  ,$      F  , ,  $T  ,$  $T  ,�  %  ,�  %  ,$  $T  ,$      F  , ,  $T  ,$  $T  ,�  %  ,�  %  ,$  $T  ,$      F  , ,  %�  ,$  %�  ,�  &�  ,�  &�  ,$  %�  ,$      F  , ,  %�  ,$  %�  ,�  &�  ,�  &�  ,$  %�  ,$      F  , ,  't  ,$  't  ,�  (<  ,�  (<  ,$  't  ,$      F  , ,  't  ,$  't  ,�  (<  ,�  (<  ,$  't  ,$      F  , ,  't  't  't  (<  (<  (<  (<  't  't  't      F  , ,  't  't  't  (<  (<  (<  (<  't  't  't      F  , ,  "�  't  "�  (<  #�  (<  #�  't  "�  't      F  , ,  "�  't  "�  (<  #�  (<  #�  't  "�  't      F  , ,  %�  %�  %�  &�  &�  &�  &�  %�  %�  %�      F  , ,  %�  %�  %�  &�  &�  &�  &�  %�  %�  %�      F  , ,  't  %�  't  &�  (<  &�  (<  %�  't  %�      F  , ,  't  %�  't  &�  (<  &�  (<  %�  't  %�      F  , ,  $T  !4  $T  !�  %  !�  %  !4  $T  !4      F  , ,  $T  !4  $T  !�  %  !�  %  !4  $T  !4      F  , ,  $T  �  $T   l  %   l  %  �  $T  �      F  , ,  $T  �  $T   l  %   l  %  �  $T  �      F  , ,  "�  "�  "�  #�  #�  #�  #�  "�  "�  "�      F  , ,  "�  "�  "�  #�  #�  #�  #�  "�  "�  "�      F  , ,  $T  "�  $T  #�  %  #�  %  "�  $T  "�      F  , ,  $T  "�  $T  #�  %  #�  %  "�  $T  "�      F  , ,  %�  "�  %�  #�  &�  #�  &�  "�  %�  "�      F  , ,  %�  "�  %�  #�  &�  #�  &�  "�  %�  "�      F  , ,  't  "�  't  #�  (<  #�  (<  "�  't  "�      F  , ,  't  "�  't  #�  (<  #�  (<  "�  't  "�      F  , ,  %�  !4  %�  !�  &�  !�  &�  !4  %�  !4      F  , ,  %�  !4  %�  !�  &�  !�  &�  !4  %�  !4      F  , ,  %�  �  %�   l  &�   l  &�  �  %�  �      F  , ,  %�  �  %�   l  &�   l  &�  �  %�  �      F  , ,  "�  !4  "�  !�  #�  !�  #�  !4  "�  !4      F  , ,  "�  !4  "�  !�  #�  !�  #�  !4  "�  !4      F  , ,  "�  $T  "�  %  #�  %  #�  $T  "�  $T      F  , ,  "�  $T  "�  %  #�  %  #�  $T  "�  $T      F  , ,  $T  $T  $T  %  %  %  %  $T  $T  $T      F  , ,  $T  $T  $T  %  %  %  %  $T  $T  $T      F  , ,  %�  $T  %�  %  &�  %  &�  $T  %�  $T      F  , ,  %�  $T  %�  %  &�  %  &�  $T  %�  $T      F  , ,  "�  �  "�   l  #�   l  #�  �  "�  �      F  , ,  "�  �  "�   l  #�   l  #�  �  "�  �      F  , ,  't  $T  't  %  (<  %  (<  $T  't  $T      F  , ,  't  $T  't  %  (<  %  (<  $T  't  $T      F  , ,  't  !4  't  !�  (<  !�  (<  !4  't  !4      F  , ,  't  !4  't  !�  (<  !�  (<  !4  't  !4      F  , ,  't  �  't   l  (<   l  (<  �  't  �      F  , ,  't  �  't   l  (<   l  (<  �  't  �      F  , ,  "�  %�  "�  &�  #�  &�  #�  %�  "�  %�      F  , ,  "�  %�  "�  &�  #�  &�  #�  %�  "�  %�      F  , ,  $T  %�  $T  &�  %  &�  %  %�  $T  %�      F  , ,  $T  %�  $T  &�  %  &�  %  %�  $T  %�      F  , ,  /D  �  /D   l  0   l  0  �  /D  �      F  , ,  /D  �  /D   l  0   l  0  �  /D  �      F  , ,  *�  "�  *�  #�  +\  #�  +\  "�  *�  "�      F  , ,  *�  "�  *�  #�  +\  #�  +\  "�  *�  "�      F  , ,  ,$  �  ,$   l  ,�   l  ,�  �  ,$  �      F  , ,  ,$  �  ,$   l  ,�   l  ,�  �  ,$  �      F  , ,  *�  $T  *�  %  +\  %  +\  $T  *�  $T      F  , ,  *�  $T  *�  %  +\  %  +\  $T  *�  $T      F  , ,  ,$  $T  ,$  %  ,�  %  ,�  $T  ,$  $T      F  , ,  ,$  $T  ,$  %  ,�  %  ,�  $T  ,$  $T      F  , ,  -�  $T  -�  %  .|  %  .|  $T  -�  $T      F  , ,  -�  $T  -�  %  .|  %  .|  $T  -�  $T      F  , ,  /D  $T  /D  %  0  %  0  $T  /D  $T      F  , ,  /D  $T  /D  %  0  %  0  $T  /D  $T      F  , ,  ,$  "�  ,$  #�  ,�  #�  ,�  "�  ,$  "�      F  , ,  ,$  "�  ,$  #�  ,�  #�  ,�  "�  ,$  "�      F  , ,  -�  "�  -�  #�  .|  #�  .|  "�  -�  "�      F  , ,  -�  "�  -�  #�  .|  #�  .|  "�  -�  "�      F  , ,  /D  "�  /D  #�  0  #�  0  "�  /D  "�      F  , ,  /D  "�  /D  #�  0  #�  0  "�  /D  "�      F  , ,  *�  �  *�   l  +\   l  +\  �  *�  �      F  , ,  *�  �  *�   l  +\   l  +\  �  *�  �      F  , ,  *�  !4  *�  !�  +\  !�  +\  !4  *�  !4      F  , ,  *�  !4  *�  !�  +\  !�  +\  !4  *�  !4      F  , ,  ,$  !4  ,$  !�  ,�  !�  ,�  !4  ,$  !4      F  , ,  ,$  !4  ,$  !�  ,�  !�  ,�  !4  ,$  !4      F  , ,  -�  �  -�   l  .|   l  .|  �  -�  �      F  , ,  -�  �  -�   l  .|   l  .|  �  -�  �      F  , ,  -�  !4  -�  !�  .|  !�  .|  !4  -�  !4      F  , ,  -�  !4  -�  !�  .|  !�  .|  !4  -�  !4      F  , ,  *�  %�  *�  &�  +\  &�  +\  %�  *�  %�      F  , ,  *�  %�  *�  &�  +\  &�  +\  %�  *�  %�      F  , ,  ,$  %�  ,$  &�  ,�  &�  ,�  %�  ,$  %�      F  , ,  ,$  %�  ,$  &�  ,�  &�  ,�  %�  ,$  %�      F  , ,  -�  %�  -�  &�  .|  &�  .|  %�  -�  %�      F  , ,  -�  %�  -�  &�  .|  &�  .|  %�  -�  %�      F  , ,  /D  %�  /D  &�  0  &�  0  %�  /D  %�      F  , ,  /D  %�  /D  &�  0  &�  0  %�  /D  %�      F  , ,  /D  !4  /D  !�  0  !�  0  !4  /D  !4      F  , ,  /D  !4  /D  !�  0  !�  0  !4  /D  !4      F  , ,  ?  &�  ?  't  ?�  't  ?�  &�  ?  &�      F  , ,  ?  &�  ?  't  ?�  't  ?�  &�  ?  &�      F  , ,  8�  ,$  8�  ,�  9l  ,�  9l  ,$  8�  ,$      F  , ,  8�  ,$  8�  ,�  9l  ,�  9l  ,$  8�  ,$      F  , ,  :4  ,$  :4  ,�  :�  ,�  :�  ,$  :4  ,$      F  , ,  :4  ,$  :4  ,�  :�  ,�  :�  ,$  :4  ,$      F  , ,  8�  't  8�  (<  9l  (<  9l  't  8�  't      F  , ,  8�  't  8�  (<  9l  (<  9l  't  8�  't      F  , ,  :4  't  :4  (<  :�  (<  :�  't  :4  't      F  , ,  :4  't  :4  (<  :�  (<  :�  't  :4  't      F  , ,  8�  )  8�  )�  9l  )�  9l  )  8�  )      F  , ,  8�  )  8�  )�  9l  )�  9l  )  8�  )      F  , ,  :4  )  :4  )�  :�  )�  :�  )  :4  )      F  , ,  :4  )  :4  )�  :�  )�  :�  )  :4  )      F  , ,  :4  *�  :4  +\  :�  +\  :�  *�  :4  *�      F  , ,  :4  *�  :4  +\  :�  +\  :�  *�  :4  *�      F  , ,  ?  (<  ?  )  ?�  )  ?�  (<  ?  (<      F  , ,  ?  (<  ?  )  ?�  )  ?�  (<  ?  (<      F  , ,  ?  )�  ?  *�  ?�  *�  ?�  )�  ?  )�      F  , ,  ?  )�  ?  *�  ?�  *�  ?�  )�  ?  )�      F  , ,  ?  +\  ?  ,$  ?�  ,$  ?�  +\  ?  +\      F  , ,  ?  +\  ?  ,$  ?�  ,$  ?�  +\  ?  +\      F  , ,  ?  ,�  ?  -�  ?�  -�  ?�  ,�  ?  ,�      F  , ,  ?  ,�  ?  -�  ?�  -�  ?�  ,�  ?  ,�      F  , ,  8�  *�  8�  +\  9l  +\  9l  *�  8�  *�      F  , ,  8�  *�  8�  +\  9l  +\  9l  *�  8�  *�      F  , ,  0�  ,$  0�  ,�  1�  ,�  1�  ,$  0�  ,$      F  , ,  0�  ,$  0�  ,�  1�  ,�  1�  ,$  0�  ,$      F  , ,  2d  ,$  2d  ,�  3,  ,�  3,  ,$  2d  ,$      F  , ,  2d  ,$  2d  ,�  3,  ,�  3,  ,$  2d  ,$      F  , ,  0�  )  0�  )�  1�  )�  1�  )  0�  )      F  , ,  0�  )  0�  )�  1�  )�  1�  )  0�  )      F  , ,  2d  )  2d  )�  3,  )�  3,  )  2d  )      F  , ,  2d  )  2d  )�  3,  )�  3,  )  2d  )      F  , ,  3�  )  3�  )�  4�  )�  4�  )  3�  )      F  , ,  3�  )  3�  )�  4�  )�  4�  )  3�  )      F  , ,  5�  )  5�  )�  6L  )�  6L  )  5�  )      F  , ,  5�  )  5�  )�  6L  )�  6L  )  5�  )      F  , ,  7  )  7  )�  7�  )�  7�  )  7  )      F  , ,  7  )  7  )�  7�  )�  7�  )  7  )      F  , ,  3�  ,$  3�  ,�  4�  ,�  4�  ,$  3�  ,$      F  , ,  3�  ,$  3�  ,�  4�  ,�  4�  ,$  3�  ,$      F  , ,  5�  ,$  5�  ,�  6L  ,�  6L  ,$  5�  ,$      F  , ,  5�  ,$  5�  ,�  6L  ,�  6L  ,$  5�  ,$      F  , ,  7  ,$  7  ,�  7�  ,�  7�  ,$  7  ,$      F  , ,  7  ,$  7  ,�  7�  ,�  7�  ,$  7  ,$      F  , ,  0�  't  0�  (<  1�  (<  1�  't  0�  't      F  , ,  0�  't  0�  (<  1�  (<  1�  't  0�  't      F  , ,  2d  't  2d  (<  3,  (<  3,  't  2d  't      F  , ,  2d  't  2d  (<  3,  (<  3,  't  2d  't      F  , ,  3�  't  3�  (<  4�  (<  4�  't  3�  't      F  , ,  3�  't  3�  (<  4�  (<  4�  't  3�  't      F  , ,  5�  't  5�  (<  6L  (<  6L  't  5�  't      F  , ,  5�  't  5�  (<  6L  (<  6L  't  5�  't      F  , ,  0�  *�  0�  +\  1�  +\  1�  *�  0�  *�      F  , ,  0�  *�  0�  +\  1�  +\  1�  *�  0�  *�      F  , ,  2d  *�  2d  +\  3,  +\  3,  *�  2d  *�      F  , ,  2d  *�  2d  +\  3,  +\  3,  *�  2d  *�      F  , ,  3�  *�  3�  +\  4�  +\  4�  *�  3�  *�      F  , ,  3�  *�  3�  +\  4�  +\  4�  *�  3�  *�      F  , ,  5�  *�  5�  +\  6L  +\  6L  *�  5�  *�      F  , ,  5�  *�  5�  +\  6L  +\  6L  *�  5�  *�      F  , ,  7  *�  7  +\  7�  +\  7�  *�  7  *�      F  , ,  7  *�  7  +\  7�  +\  7�  *�  7  *�      F  , ,  7  't  7  (<  7�  (<  7�  't  7  't      F  , ,  7  't  7  (<  7�  (<  7�  't  7  't      F  , ,  3�  �  3�   l  4�   l  4�  �  3�  �      F  , ,  3�  �  3�   l  4�   l  4�  �  3�  �      F  , ,  0�  $T  0�  %  1�  %  1�  $T  0�  $T      F  , ,  0�  $T  0�  %  1�  %  1�  $T  0�  $T      F  , ,  2d  $T  2d  %  3,  %  3,  $T  2d  $T      F  , ,  2d  $T  2d  %  3,  %  3,  $T  2d  $T      F  , ,  3�  $T  3�  %  4�  %  4�  $T  3�  $T      F  , ,  3�  $T  3�  %  4�  %  4�  $T  3�  $T      F  , ,  2d  !4  2d  !�  3,  !�  3,  !4  2d  !4      F  , ,  2d  !4  2d  !�  3,  !�  3,  !4  2d  !4      F  , ,  0�  %�  0�  &�  1�  &�  1�  %�  0�  %�      F  , ,  0�  %�  0�  &�  1�  &�  1�  %�  0�  %�      F  , ,  7  �  7   l  7�   l  7�  �  7  �      F  , ,  7  �  7   l  7�   l  7�  �  7  �      F  , ,  2d  %�  2d  &�  3,  &�  3,  %�  2d  %�      F  , ,  2d  %�  2d  &�  3,  &�  3,  %�  2d  %�      F  , ,  3�  %�  3�  &�  4�  &�  4�  %�  3�  %�      F  , ,  3�  %�  3�  &�  4�  &�  4�  %�  3�  %�      F  , ,  5�  %�  5�  &�  6L  &�  6L  %�  5�  %�      F  , ,  5�  %�  5�  &�  6L  &�  6L  %�  5�  %�      F  , ,  7  %�  7  &�  7�  &�  7�  %�  7  %�      F  , ,  7  %�  7  &�  7�  &�  7�  %�  7  %�      F  , ,  5�  $T  5�  %  6L  %  6L  $T  5�  $T      F  , ,  5�  $T  5�  %  6L  %  6L  $T  5�  $T      F  , ,  5�  "�  5�  #�  6L  #�  6L  "�  5�  "�      F  , ,  5�  "�  5�  #�  6L  #�  6L  "�  5�  "�      F  , ,  7  "�  7  #�  7�  #�  7�  "�  7  "�      F  , ,  7  "�  7  #�  7�  #�  7�  "�  7  "�      F  , ,  5�  �  5�   l  6L   l  6L  �  5�  �      F  , ,  5�  �  5�   l  6L   l  6L  �  5�  �      F  , ,  5�  !4  5�  !�  6L  !�  6L  !4  5�  !4      F  , ,  5�  !4  5�  !�  6L  !�  6L  !4  5�  !4      F  , ,  3�  !4  3�  !�  4�  !�  4�  !4  3�  !4      F  , ,  3�  !4  3�  !�  4�  !�  4�  !4  3�  !4      F  , ,  0�  "�  0�  #�  1�  #�  1�  "�  0�  "�      F  , ,  0�  "�  0�  #�  1�  #�  1�  "�  0�  "�      F  , ,  7  !4  7  !�  7�  !�  7�  !4  7  !4      F  , ,  7  !4  7  !�  7�  !�  7�  !4  7  !4      F  , ,  2d  �  2d   l  3,   l  3,  �  2d  �      F  , ,  2d  �  2d   l  3,   l  3,  �  2d  �      F  , ,  0�  !4  0�  !�  1�  !�  1�  !4  0�  !4      F  , ,  0�  !4  0�  !�  1�  !�  1�  !4  0�  !4      F  , ,  7  $T  7  %  7�  %  7�  $T  7  $T      F  , ,  7  $T  7  %  7�  %  7�  $T  7  $T      F  , ,  2d  "�  2d  #�  3,  #�  3,  "�  2d  "�      F  , ,  2d  "�  2d  #�  3,  #�  3,  "�  2d  "�      F  , ,  0�  �  0�   l  1�   l  1�  �  0�  �      F  , ,  0�  �  0�   l  1�   l  1�  �  0�  �      F  , ,  3�  "�  3�  #�  4�  #�  4�  "�  3�  "�      F  , ,  3�  "�  3�  #�  4�  #�  4�  "�  3�  "�      F  , ,  8�  "�  8�  #�  9l  #�  9l  "�  8�  "�      F  , ,  8�  "�  8�  #�  9l  #�  9l  "�  8�  "�      F  , ,  8�  �  8�   l  9l   l  9l  �  8�  �      F  , ,  8�  �  8�   l  9l   l  9l  �  8�  �      F  , ,  :4  "�  :4  #�  :�  #�  :�  "�  :4  "�      F  , ,  :4  "�  :4  #�  :�  #�  :�  "�  :4  "�      F  , ,  :4  $T  :4  %  :�  %  :�  $T  :4  $T      F  , ,  :4  $T  :4  %  :�  %  :�  $T  :4  $T      F  , ,  :4  %�  :4  &�  :�  &�  :�  %�  :4  %�      F  , ,  :4  %�  :4  &�  :�  &�  :�  %�  :4  %�      F  , ,  8�  $T  8�  %  9l  %  9l  $T  8�  $T      F  , ,  8�  $T  8�  %  9l  %  9l  $T  8�  $T      F  , ,  8�  !4  8�  !�  9l  !�  9l  !4  8�  !4      F  , ,  8�  !4  8�  !�  9l  !�  9l  !4  8�  !4      F  , ,  :4  !4  :4  !�  :�  !�  :�  !4  :4  !4      F  , ,  :4  !4  :4  !�  :�  !�  :�  !4  :4  !4      F  , ,  8�  %�  8�  &�  9l  &�  9l  %�  8�  %�      F  , ,  8�  %�  8�  &�  9l  &�  9l  %�  8�  %�      F  , ,  ?   l  ?  !4  ?�  !4  ?�   l  ?   l      F  , ,  ?   l  ?  !4  ?�  !4  ?�   l  ?   l      F  , ,  ?  !�  ?  "�  ?�  "�  ?�  !�  ?  !�      F  , ,  ?  !�  ?  "�  ?�  "�  ?�  !�  ?  !�      F  , ,  ?  #�  ?  $T  ?�  $T  ?�  #�  ?  #�      F  , ,  ?  #�  ?  $T  ?�  $T  ?�  #�  ?  #�      F  , ,  ?  %  ?  %�  ?�  %�  ?�  %  ?  %      F  , ,  ?  %  ?  %�  ?�  %�  ?�  %  ?  %      F  , ,  :4  �  :4   l  :�   l  :�  �  :4  �      F  , ,  :4  �  :4   l  :�   l  :�  �  :4  �      F  , ,  �  -�  �  .|  l  .|  l  -�  �  -�      F  , ,  �  -�  �  .|  l  .|  l  -�  �  -�      F  , ,  4  -�  4  .|  �  .|  �  -�  4  -�      F  , ,  4  -�  4  .|  �  .|  �  -�  4  -�      F  , ,  	�  -�  	�  .|  
�  .|  
�  -�  	�  -�      F  , ,  	�  -�  	�  .|  
�  .|  
�  -�  	�  -�      F  , ,  T  -�  T  .|    .|    -�  T  -�      F  , ,  T  -�  T  .|    .|    -�  T  -�      F  , ,  �  -�  �  .|  �  .|  �  -�  �  -�      F  , ,  �  -�  �  .|  �  .|  �  -�  �  -�      F  , ,  t  -�  t  .|  <  .|  <  -�  t  -�      F  , ,  t  -�  t  .|  <  .|  <  -�  t  -�      F  , ,    -�    .|  �  .|  �  -�    -�      F  , ,    -�    .|  �  .|  �  -�    -�      F  , ,  �  -�  �  .|  \  .|  \  -�  �  -�      F  , ,  �  -�  �  .|  \  .|  \  -�  �  -�      F  , ,  $  -�  $  .|  �  .|  �  -�  $  -�      F  , ,  $  -�  $  .|  �  .|  �  -�  $  -�      F  , ,  �  -�  �  .|  |  .|  |  -�  �  -�      F  , ,  �  -�  �  .|  |  .|  |  -�  �  -�      F  , ,  D  -�  D  .|    .|    -�  D  -�      F  , ,  D  -�  D  .|    .|    -�  D  -�      F  , ,  �  -�  �  .|  �  .|  �  -�  �  -�      F  , ,  �  -�  �  .|  �  .|  �  -�  �  -�      F  , ,  d  -�  d  .|  ,  .|  ,  -�  d  -�      F  , ,  d  -�  d  .|  ,  .|  ,  -�  d  -�      F  , ,  �  -�  �  .|  �  .|  �  -�  �  -�      F  , ,  �  -�  �  .|  �  .|  �  -�  �  -�      F  , ,  �  -�  �  .|  L  .|  L  -�  �  -�      F  , ,  �  -�  �  .|  L  .|  L  -�  �  -�      F  , ,    -�    .|  �  .|  �  -�    -�      F  , ,    -�    .|  �  .|  �  -�    -�      F  , ,  �  -�  �  .|   l  .|   l  -�  �  -�      F  , ,  �  -�  �  .|   l  .|   l  -�  �  -�      F  , ,  �  -�  �  .|  L  .|  L  -�  �  -�      F  , ,  �  -�  �  .|  L  .|  L  -�  �  -�      F  , ,    -�    .|  �  .|  �  -�    -�      F  , ,    -�    .|  �  .|  �  -�    -�      F  , ,  d  /D  d  0  ,  0  ,  /D  d  /D      F  , ,  d  /D  d  0  ,  0  ,  /D  d  /D      F  , ,  d  0�  d  1�  ,  1�  ,  0�  d  0�      F  , ,  d  0�  d  1�  ,  1�  ,  0�  d  0�      F  , ,  d  2d  d  3,  ,  3,  ,  2d  d  2d      F  , ,  d  2d  d  3,  ,  3,  ,  2d  d  2d      F  , ,  d  3�  d  4�  ,  4�  ,  3�  d  3�      F  , ,  d  3�  d  4�  ,  4�  ,  3�  d  3�      F  , ,  $  5�  $  6L  �  6L  �  5�  $  5�      F  , ,  $  5�  $  6L  �  6L  �  5�  $  5�      F  , ,  �  5�  �  6L  |  6L  |  5�  �  5�      F  , ,  �  5�  �  6L  |  6L  |  5�  �  5�      F  , ,  D  5�  D  6L    6L    5�  D  5�      F  , ,  D  5�  D  6L    6L    5�  D  5�      F  , ,  �  5�  �  6L  �  6L  �  5�  �  5�      F  , ,  �  5�  �  6L  �  6L  �  5�  �  5�      F  , ,  d  5�  d  6L  ,  6L  ,  5�  d  5�      F  , ,  d  5�  d  6L  ,  6L  ,  5�  d  5�      F  , ,  �  5�  �  6L  �  6L  �  5�  �  5�      F  , ,  �  5�  �  6L  �  6L  �  5�  �  5�      F  , ,  �  5�  �  6L  L  6L  L  5�  �  5�      F  , ,  �  5�  �  6L  L  6L  L  5�  �  5�      F  , ,    5�    6L  �  6L  �  5�    5�      F  , ,    5�    6L  �  6L  �  5�    5�      F  , ,  �  5�  �  6L   l  6L   l  5�  �  5�      F  , ,  �  5�  �  6L   l  6L   l  5�  �  5�      F  , ,  d  7  d  7�  ,  7�  ,  7  d  7      F  , ,  d  7  d  7�  ,  7�  ,  7  d  7      F  , ,  d  8�  d  9l  ,  9l  ,  8�  d  8�      F  , ,  d  8�  d  9l  ,  9l  ,  8�  d  8�      F  , ,  d  :4  d  :�  ,  :�  ,  :4  d  :4      F  , ,  d  :4  d  :�  ,  :�  ,  :4  d  :4      F  , ,    7    7�  �  7�  �  7    7      F  , ,    7    7�  �  7�  �  7    7      F  , ,  �  7  �  7�   l  7�   l  7  �  7      F  , ,  �  7  �  7�   l  7�   l  7  �  7      F  , ,  �  7  �  7�  �  7�  �  7  �  7      F  , ,  �  7  �  7�  �  7�  �  7  �  7      F  , ,  �  8�  �  9l  �  9l  �  8�  �  8�      F  , ,  �  8�  �  9l  �  9l  �  8�  �  8�      F  , ,  �  8�  �  9l  L  9l  L  8�  �  8�      F  , ,  �  8�  �  9l  L  9l  L  8�  �  8�      F  , ,    8�    9l  �  9l  �  8�    8�      F  , ,    8�    9l  �  9l  �  8�    8�      F  , ,  �  8�  �  9l   l  9l   l  8�  �  8�      F  , ,  �  8�  �  9l   l  9l   l  8�  �  8�      F  , ,  �  7  �  7�  L  7�  L  7  �  7      F  , ,  �  7  �  7�  L  7�  L  7  �  7      F  , ,  �  :4  �  :�  �  :�  �  :4  �  :4      F  , ,  �  :4  �  :�  �  :�  �  :4  �  :4      F  , ,  �  :4  �  :�  L  :�  L  :4  �  :4      F  , ,  �  :4  �  :�  L  :�  L  :4  �  :4      F  , ,    :4    :�  �  :�  �  :4    :4      F  , ,    :4    :�  �  :�  �  :4    :4      F  , ,  �  :4  �  :�   l  :�   l  :4  �  :4      F  , ,  �  :4  �  :�   l  :�   l  :4  �  :4      F  , ,  �  7  �  7�  �  7�  �  7  �  7      F  , ,  �  7  �  7�  �  7�  �  7  �  7      F  , ,  $  7  $  7�  �  7�  �  7  $  7      F  , ,  $  7  $  7�  �  7�  �  7  $  7      F  , ,  $  8�  $  9l  �  9l  �  8�  $  8�      F  , ,  $  8�  $  9l  �  9l  �  8�  $  8�      F  , ,  $  :4  $  :�  �  :�  �  :4  $  :4      F  , ,  $  :4  $  :�  �  :�  �  :4  $  :4      F  , ,  �  :4  �  :�  |  :�  |  :4  �  :4      F  , ,  �  :4  �  :�  |  :�  |  :4  �  :4      F  , ,  D  :4  D  :�    :�    :4  D  :4      F  , ,  D  :4  D  :�    :�    :4  D  :4      F  , ,  �  :4  �  :�  �  :�  �  :4  �  :4      F  , ,  �  :4  �  :�  �  :�  �  :4  �  :4      F  , ,  �  8�  �  9l  |  9l  |  8�  �  8�      F  , ,  �  8�  �  9l  |  9l  |  8�  �  8�      F  , ,  D  8�  D  9l    9l    8�  D  8�      F  , ,  D  8�  D  9l    9l    8�  D  8�      F  , ,  �  8�  �  9l  �  9l  �  8�  �  8�      F  , ,  �  8�  �  9l  �  9l  �  8�  �  8�      F  , ,  �  7  �  7�  |  7�  |  7  �  7      F  , ,  �  7  �  7�  |  7�  |  7  �  7      F  , ,  D  7  D  7�    7�    7  D  7      F  , ,  D  7  D  7�    7�    7  D  7      F  , ,  D  /D  D  0    0    /D  D  /D      F  , ,  D  /D  D  0    0    /D  D  /D      F  , ,  $  3�  $  4�  �  4�  �  3�  $  3�      F  , ,  $  3�  $  4�  �  4�  �  3�  $  3�      F  , ,  �  3�  �  4�  |  4�  |  3�  �  3�      F  , ,  �  3�  �  4�  |  4�  |  3�  �  3�      F  , ,  D  3�  D  4�    4�    3�  D  3�      F  , ,  D  3�  D  4�    4�    3�  D  3�      F  , ,  �  3�  �  4�  �  4�  �  3�  �  3�      F  , ,  �  3�  �  4�  �  4�  �  3�  �  3�      F  , ,  $  0�  $  1�  �  1�  �  0�  $  0�      F  , ,  $  0�  $  1�  �  1�  �  0�  $  0�      F  , ,  �  0�  �  1�  |  1�  |  0�  �  0�      F  , ,  �  0�  �  1�  |  1�  |  0�  �  0�      F  , ,  D  0�  D  1�    1�    0�  D  0�      F  , ,  D  0�  D  1�    1�    0�  D  0�      F  , ,  �  0�  �  1�  �  1�  �  0�  �  0�      F  , ,  �  0�  �  1�  �  1�  �  0�  �  0�      F  , ,  �  /D  �  0  �  0  �  /D  �  /D      F  , ,  �  /D  �  0  �  0  �  /D  �  /D      F  , ,  $  2d  $  3,  �  3,  �  2d  $  2d      F  , ,  $  2d  $  3,  �  3,  �  2d  $  2d      F  , ,  �  2d  �  3,  |  3,  |  2d  �  2d      F  , ,  �  2d  �  3,  |  3,  |  2d  �  2d      F  , ,  D  2d  D  3,    3,    2d  D  2d      F  , ,  D  2d  D  3,    3,    2d  D  2d      F  , ,  �  2d  �  3,  �  3,  �  2d  �  2d      F  , ,  �  2d  �  3,  �  3,  �  2d  �  2d      F  , ,  $  /D  $  0  �  0  �  /D  $  /D      F  , ,  $  /D  $  0  �  0  �  /D  $  /D      F  , ,  �  /D  �  0  |  0  |  /D  �  /D      F  , ,  �  /D  �  0  |  0  |  /D  �  /D      F  , ,  �  2d  �  3,   l  3,   l  2d  �  2d      F  , ,  �  2d  �  3,   l  3,   l  2d  �  2d      F  , ,  �  0�  �  1�  L  1�  L  0�  �  0�      F  , ,  �  0�  �  1�  L  1�  L  0�  �  0�      F  , ,    0�    1�  �  1�  �  0�    0�      F  , ,    0�    1�  �  1�  �  0�    0�      F  , ,  �  0�  �  1�   l  1�   l  0�  �  0�      F  , ,  �  0�  �  1�   l  1�   l  0�  �  0�      F  , ,  �  /D  �  0  L  0  L  /D  �  /D      F  , ,  �  /D  �  0  L  0  L  /D  �  /D      F  , ,    /D    0  �  0  �  /D    /D      F  , ,    /D    0  �  0  �  /D    /D      F  , ,  �  3�  �  4�  �  4�  �  3�  �  3�      F  , ,  �  3�  �  4�  �  4�  �  3�  �  3�      F  , ,  �  3�  �  4�  L  4�  L  3�  �  3�      F  , ,  �  3�  �  4�  L  4�  L  3�  �  3�      F  , ,    3�    4�  �  4�  �  3�    3�      F  , ,    3�    4�  �  4�  �  3�    3�      F  , ,  �  3�  �  4�   l  4�   l  3�  �  3�      F  , ,  �  3�  �  4�   l  4�   l  3�  �  3�      F  , ,  �  /D  �  0   l  0   l  /D  �  /D      F  , ,  �  /D  �  0   l  0   l  /D  �  /D      F  , ,  �  /D  �  0  �  0  �  /D  �  /D      F  , ,  �  /D  �  0  �  0  �  /D  �  /D      F  , ,  �  0�  �  1�  �  1�  �  0�  �  0�      F  , ,  �  0�  �  1�  �  1�  �  0�  �  0�      F  , ,  �  2d  �  3,  �  3,  �  2d  �  2d      F  , ,  �  2d  �  3,  �  3,  �  2d  �  2d      F  , ,  �  2d  �  3,  L  3,  L  2d  �  2d      F  , ,  �  2d  �  3,  L  3,  L  2d  �  2d      F  , ,    2d    3,  �  3,  �  2d    2d      F  , ,    2d    3,  �  3,  �  2d    2d      F  , ,  �  5�  �  6L  L  6L  L  5�  �  5�      F  , ,  �  5�  �  6L  L  6L  L  5�  �  5�      F  , ,    5�    6L  �  6L  �  5�    5�      F  , ,    5�    6L  �  6L  �  5�    5�      F  , ,  �  5�  �  6L  l  6L  l  5�  �  5�      F  , ,  �  5�  �  6L  l  6L  l  5�  �  5�      F  , ,  4  5�  4  6L  �  6L  �  5�  4  5�      F  , ,  4  5�  4  6L  �  6L  �  5�  4  5�      F  , ,  	�  5�  	�  6L  
�  6L  
�  5�  	�  5�      F  , ,  	�  5�  	�  6L  
�  6L  
�  5�  	�  5�      F  , ,  T  5�  T  6L    6L    5�  T  5�      F  , ,  T  5�  T  6L    6L    5�  T  5�      F  , ,  �  5�  �  6L  �  6L  �  5�  �  5�      F  , ,  �  5�  �  6L  �  6L  �  5�  �  5�      F  , ,  t  5�  t  6L  <  6L  <  5�  t  5�      F  , ,  t  5�  t  6L  <  6L  <  5�  t  5�      F  , ,    5�    6L  �  6L  �  5�    5�      F  , ,    5�    6L  �  6L  �  5�    5�      F  , ,  �  5�  �  6L  \  6L  \  5�  �  5�      F  , ,  �  5�  �  6L  \  6L  \  5�  �  5�      F  , ,  T  7  T  7�    7�    7  T  7      F  , ,  T  7  T  7�    7�    7  T  7      F  , ,  �  7  �  7�  �  7�  �  7  �  7      F  , ,  �  7  �  7�  �  7�  �  7  �  7      F  , ,  t  7  t  7�  <  7�  <  7  t  7      F  , ,  t  7  t  7�  <  7�  <  7  t  7      F  , ,    7    7�  �  7�  �  7    7      F  , ,    7    7�  �  7�  �  7    7      F  , ,  �  7  �  7�  \  7�  \  7  �  7      F  , ,  �  7  �  7�  \  7�  \  7  �  7      F  , ,  T  8�  T  9l    9l    8�  T  8�      F  , ,  T  8�  T  9l    9l    8�  T  8�      F  , ,  �  8�  �  9l  �  9l  �  8�  �  8�      F  , ,  �  8�  �  9l  �  9l  �  8�  �  8�      F  , ,  t  8�  t  9l  <  9l  <  8�  t  8�      F  , ,  t  8�  t  9l  <  9l  <  8�  t  8�      F  , ,    8�    9l  �  9l  �  8�    8�      F  , ,    8�    9l  �  9l  �  8�    8�      F  , ,  �  8�  �  9l  \  9l  \  8�  �  8�      F  , ,  �  8�  �  9l  \  9l  \  8�  �  8�      F  , ,  T  :4  T  :�    :�    :4  T  :4      F  , ,  T  :4  T  :�    :�    :4  T  :4      F  , ,  �  :4  �  :�  �  :�  �  :4  �  :4      F  , ,  �  :4  �  :�  �  :�  �  :4  �  :4      F  , ,  t  :4  t  :�  <  :�  <  :4  t  :4      F  , ,  t  :4  t  :�  <  :�  <  :4  t  :4      F  , ,    :4    :�  �  :�  �  :4    :4      F  , ,    :4    :�  �  :�  �  :4    :4      F  , ,  �  :4  �  :�  \  :�  \  :4  �  :4      F  , ,  �  :4  �  :�  \  :�  \  :4  �  :4      F  , ,  �  7  �  7�  L  7�  L  7  �  7      F  , ,  �  7  �  7�  L  7�  L  7  �  7      F  , ,    7    7�  �  7�  �  7    7      F  , ,    7    7�  �  7�  �  7    7      F  , ,  �  7  �  7�  l  7�  l  7  �  7      F  , ,  �  7  �  7�  l  7�  l  7  �  7      F  , ,  4  7  4  7�  �  7�  �  7  4  7      F  , ,  4  7  4  7�  �  7�  �  7  4  7      F  , ,  	�  7  	�  7�  
�  7�  
�  7  	�  7      F  , ,  	�  7  	�  7�  
�  7�  
�  7  	�  7      F  , ,  �  :4  �  :�  L  :�  L  :4  �  :4      F  , ,  �  :4  �  :�  L  :�  L  :4  �  :4      F  , ,    :4    :�  �  :�  �  :4    :4      F  , ,    :4    :�  �  :�  �  :4    :4      F  , ,  �  :4  �  :�  l  :�  l  :4  �  :4      F  , ,  �  :4  �  :�  l  :�  l  :4  �  :4      F  , ,  4  :4  4  :�  �  :�  �  :4  4  :4      F  , ,  4  :4  4  :�  �  :�  �  :4  4  :4      F  , ,  	�  :4  	�  :�  
�  :�  
�  :4  	�  :4      F  , ,  	�  :4  	�  :�  
�  :�  
�  :4  	�  :4      F  , ,  �  8�  �  9l  L  9l  L  8�  �  8�      F  , ,  �  8�  �  9l  L  9l  L  8�  �  8�      F  , ,    8�    9l  �  9l  �  8�    8�      F  , ,    8�    9l  �  9l  �  8�    8�      F  , ,  �  8�  �  9l  l  9l  l  8�  �  8�      F  , ,  �  8�  �  9l  l  9l  l  8�  �  8�      F  , ,  4  8�  4  9l  �  9l  �  8�  4  8�      F  , ,  4  8�  4  9l  �  9l  �  8�  4  8�      F  , ,  	�  8�  	�  9l  
�  9l  
�  8�  	�  8�      F  , ,  	�  8�  	�  9l  
�  9l  
�  8�  	�  8�      F  , ,  4  0�  4  1�  �  1�  �  0�  4  0�      F  , ,  4  0�  4  1�  �  1�  �  0�  4  0�      F  , ,  �  3�  �  4�  L  4�  L  3�  �  3�      F  , ,  �  3�  �  4�  L  4�  L  3�  �  3�      F  , ,    3�    4�  �  4�  �  3�    3�      F  , ,    3�    4�  �  4�  �  3�    3�      F  , ,  �  3�  �  4�  l  4�  l  3�  �  3�      F  , ,  �  3�  �  4�  l  4�  l  3�  �  3�      F  , ,  4  3�  4  4�  �  4�  �  3�  4  3�      F  , ,  4  3�  4  4�  �  4�  �  3�  4  3�      F  , ,  	�  3�  	�  4�  
�  4�  
�  3�  	�  3�      F  , ,  	�  3�  	�  4�  
�  4�  
�  3�  	�  3�      F  , ,  	�  0�  	�  1�  
�  1�  
�  0�  	�  0�      F  , ,  	�  0�  	�  1�  
�  1�  
�  0�  	�  0�      F  , ,  4  2d  4  3,  �  3,  �  2d  4  2d      F  , ,  4  2d  4  3,  �  3,  �  2d  4  2d      F  , ,  	�  2d  	�  3,  
�  3,  
�  2d  	�  2d      F  , ,  	�  2d  	�  3,  
�  3,  
�  2d  	�  2d      F  , ,  	�  /D  	�  0  
�  0  
�  /D  	�  /D      F  , ,  	�  /D  	�  0  
�  0  
�  /D  	�  /D      F  , ,  �  2d  �  3,  L  3,  L  2d  �  2d      F  , ,  �  2d  �  3,  L  3,  L  2d  �  2d      F  , ,    2d    3,  �  3,  �  2d    2d      F  , ,    2d    3,  �  3,  �  2d    2d      F  , ,  �  2d  �  3,  l  3,  l  2d  �  2d      F  , ,  �  2d  �  3,  l  3,  l  2d  �  2d      F  , ,  �  0�  �  1�  L  1�  L  0�  �  0�      F  , ,  �  0�  �  1�  L  1�  L  0�  �  0�      F  , ,    0�    1�  �  1�  �  0�    0�      F  , ,    0�    1�  �  1�  �  0�    0�      F  , ,  �  0�  �  1�  l  1�  l  0�  �  0�      F  , ,  �  0�  �  1�  l  1�  l  0�  �  0�      F  , ,  �  /D  �  0  L  0  L  /D  �  /D      F  , ,  �  /D  �  0  L  0  L  /D  �  /D      F  , ,    /D    0  �  0  �  /D    /D      F  , ,    /D    0  �  0  �  /D    /D      F  , ,  �  /D  �  0  l  0  l  /D  �  /D      F  , ,  �  /D  �  0  l  0  l  /D  �  /D      F  , ,  4  /D  4  0  �  0  �  /D  4  /D      F  , ,  4  /D  4  0  �  0  �  /D  4  /D      F  , ,  T  2d  T  3,    3,    2d  T  2d      F  , ,  T  2d  T  3,    3,    2d  T  2d      F  , ,  �  2d  �  3,  �  3,  �  2d  �  2d      F  , ,  �  2d  �  3,  �  3,  �  2d  �  2d      F  , ,  t  2d  t  3,  <  3,  <  2d  t  2d      F  , ,  t  2d  t  3,  <  3,  <  2d  t  2d      F  , ,  T  0�  T  1�    1�    0�  T  0�      F  , ,  T  0�  T  1�    1�    0�  T  0�      F  , ,  �  0�  �  1�  �  1�  �  0�  �  0�      F  , ,  �  0�  �  1�  �  1�  �  0�  �  0�      F  , ,  t  0�  t  1�  <  1�  <  0�  t  0�      F  , ,  t  0�  t  1�  <  1�  <  0�  t  0�      F  , ,    2d    3,  �  3,  �  2d    2d      F  , ,    2d    3,  �  3,  �  2d    2d      F  , ,  �  2d  �  3,  \  3,  \  2d  �  2d      F  , ,  �  2d  �  3,  \  3,  \  2d  �  2d      F  , ,    /D    0  �  0  �  /D    /D      F  , ,    /D    0  �  0  �  /D    /D      F  , ,  �  3�  �  4�  �  4�  �  3�  �  3�      F  , ,  �  3�  �  4�  �  4�  �  3�  �  3�      F  , ,  t  3�  t  4�  <  4�  <  3�  t  3�      F  , ,  t  3�  t  4�  <  4�  <  3�  t  3�      F  , ,    3�    4�  �  4�  �  3�    3�      F  , ,    3�    4�  �  4�  �  3�    3�      F  , ,  �  3�  �  4�  \  4�  \  3�  �  3�      F  , ,  �  3�  �  4�  \  4�  \  3�  �  3�      F  , ,    0�    1�  �  1�  �  0�    0�      F  , ,    0�    1�  �  1�  �  0�    0�      F  , ,  �  0�  �  1�  \  1�  \  0�  �  0�      F  , ,  �  0�  �  1�  \  1�  \  0�  �  0�      F  , ,  �  /D  �  0  \  0  \  /D  �  /D      F  , ,  �  /D  �  0  \  0  \  /D  �  /D      F  , ,  t  /D  t  0  <  0  <  /D  t  /D      F  , ,  t  /D  t  0  <  0  <  /D  t  /D      F  , ,  T  /D  T  0    0    /D  T  /D      F  , ,  T  /D  T  0    0    /D  T  /D      F  , ,  T  3�  T  4�    4�    3�  T  3�      F  , ,  T  3�  T  4�    4�    3�  T  3�      F  , ,  �  /D  �  0  �  0  �  /D  �  /D      F  , ,  �  /D  �  0  �  0  �  /D  �  /D      F  , ,  T  't  T  (<    (<    't  T  't      F  , ,  T  't  T  (<    (<    't  T  't      F  , ,  �  't  �  (<  �  (<  �  't  �  't      F  , ,  �  't  �  (<  �  (<  �  't  �  't      F  , ,  T  )  T  )�    )�    )  T  )      F  , ,  T  )  T  )�    )�    )  T  )      F  , ,  �  )  �  )�  �  )�  �  )  �  )      F  , ,  �  )  �  )�  �  )�  �  )  �  )      F  , ,  t  )  t  )�  <  )�  <  )  t  )      F  , ,  t  )  t  )�  <  )�  <  )  t  )      F  , ,  T  *�  T  +\    +\    *�  T  *�      F  , ,  T  *�  T  +\    +\    *�  T  *�      F  , ,  �  *�  �  +\  �  +\  �  *�  �  *�      F  , ,  �  *�  �  +\  �  +\  �  *�  �  *�      F  , ,  t  *�  t  +\  <  +\  <  *�  t  *�      F  , ,  t  *�  t  +\  <  +\  <  *�  t  *�      F  , ,    *�    +\  �  +\  �  *�    *�      F  , ,    *�    +\  �  +\  �  *�    *�      F  , ,  �  *�  �  +\  \  +\  \  *�  �  *�      F  , ,  �  *�  �  +\  \  +\  \  *�  �  *�      F  , ,    )    )�  �  )�  �  )    )      F  , ,    )    )�  �  )�  �  )    )      F  , ,  �  )  �  )�  \  )�  \  )  �  )      F  , ,  �  )  �  )�  \  )�  \  )  �  )      F  , ,  t  't  t  (<  <  (<  <  't  t  't      F  , ,  t  't  t  (<  <  (<  <  't  t  't      F  , ,    't    (<  �  (<  �  't    't      F  , ,    't    (<  �  (<  �  't    't      F  , ,  �  't  �  (<  \  (<  \  't  �  't      F  , ,  �  't  �  (<  \  (<  \  't  �  't      F  , ,  T  ,$  T  ,�    ,�    ,$  T  ,$      F  , ,  T  ,$  T  ,�    ,�    ,$  T  ,$      F  , ,  �  ,$  �  ,�  �  ,�  �  ,$  �  ,$      F  , ,  �  ,$  �  ,�  �  ,�  �  ,$  �  ,$      F  , ,  t  ,$  t  ,�  <  ,�  <  ,$  t  ,$      F  , ,  t  ,$  t  ,�  <  ,�  <  ,$  t  ,$      F  , ,    ,$    ,�  �  ,�  �  ,$    ,$      F  , ,    ,$    ,�  �  ,�  �  ,$    ,$      F  , ,  �  ,$  �  ,�  \  ,�  \  ,$  �  ,$      F  , ,  �  ,$  �  ,�  \  ,�  \  ,$  �  ,$      F  , ,  �  )  �  )�  L  )�  L  )  �  )      F  , ,  �  )  �  )�  L  )�  L  )  �  )      F  , ,    )    )�  �  )�  �  )    )      F  , ,    )    )�  �  )�  �  )    )      F  , ,  �  )  �  )�  l  )�  l  )  �  )      F  , ,  �  )  �  )�  l  )�  l  )  �  )      F  , ,  4  )  4  )�  �  )�  �  )  4  )      F  , ,  4  )  4  )�  �  )�  �  )  4  )      F  , ,  	�  )  	�  )�  
�  )�  
�  )  	�  )      F  , ,  	�  )  	�  )�  
�  )�  
�  )  	�  )      F  , ,  �  ,$  �  ,�  L  ,�  L  ,$  �  ,$      F  , ,  �  ,$  �  ,�  L  ,�  L  ,$  �  ,$      F  , ,    't    (<  �  (<  �  't    't      F  , ,    't    (<  �  (<  �  't    't      F  , ,  �  't  �  (<  l  (<  l  't  �  't      F  , ,  �  't  �  (<  l  (<  l  't  �  't      F  , ,  �  *�  �  +\  L  +\  L  *�  �  *�      F  , ,  �  *�  �  +\  L  +\  L  *�  �  *�      F  , ,    *�    +\  �  +\  �  *�    *�      F  , ,    *�    +\  �  +\  �  *�    *�      F  , ,  �  *�  �  +\  l  +\  l  *�  �  *�      F  , ,  �  *�  �  +\  l  +\  l  *�  �  *�      F  , ,    ,$    ,�  �  ,�  �  ,$    ,$      F  , ,    ,$    ,�  �  ,�  �  ,$    ,$      F  , ,  �  ,$  �  ,�  l  ,�  l  ,$  �  ,$      F  , ,  �  ,$  �  ,�  l  ,�  l  ,$  �  ,$      F  , ,  4  ,$  4  ,�  �  ,�  �  ,$  4  ,$      F  , ,  4  ,$  4  ,�  �  ,�  �  ,$  4  ,$      F  , ,  	�  ,$  	�  ,�  
�  ,�  
�  ,$  	�  ,$      F  , ,  	�  ,$  	�  ,�  
�  ,�  
�  ,$  	�  ,$      F  , ,  4  't  4  (<  �  (<  �  't  4  't      F  , ,  4  't  4  (<  �  (<  �  't  4  't      F  , ,  	�  't  	�  (<  
�  (<  
�  't  	�  't      F  , ,  	�  't  	�  (<  
�  (<  
�  't  	�  't      F  , ,  4  *�  4  +\  �  +\  �  *�  4  *�      F  , ,  4  *�  4  +\  �  +\  �  *�  4  *�      F  , ,  	�  *�  	�  +\  
�  +\  
�  *�  	�  *�      F  , ,  	�  *�  	�  +\  
�  +\  
�  *�  	�  *�      F  , ,  �  't  �  (<  L  (<  L  't  �  't      F  , ,  �  't  �  (<  L  (<  L  't  �  't      F  , ,  4  $T  4  %  �  %  �  $T  4  $T      F  , ,  4  $T  4  %  �  %  �  $T  4  $T      F  , ,  	�  $T  	�  %  
�  %  
�  $T  	�  $T      F  , ,  	�  $T  	�  %  
�  %  
�  $T  	�  $T      F  , ,    !4    !�  �  !�  �  !4    !4      F  , ,    !4    !�  �  !�  �  !4    !4      F  , ,  �  !4  �  !�  l  !�  l  !4  �  !4      F  , ,  �  !4  �  !�  l  !�  l  !4  �  !4      F  , ,  4  !4  4  !�  �  !�  �  !4  4  !4      F  , ,  4  !4  4  !�  �  !�  �  !4  4  !4      F  , ,  �  "�  �  #�  L  #�  L  "�  �  "�      F  , ,  �  "�  �  #�  L  #�  L  "�  �  "�      F  , ,    "�    #�  �  #�  �  "�    "�      F  , ,    "�    #�  �  #�  �  "�    "�      F  , ,  4  "�  4  #�  �  #�  �  "�  4  "�      F  , ,  4  "�  4  #�  �  #�  �  "�  4  "�      F  , ,  �  �  �   l  L   l  L  �  �  �      F  , ,  �  �  �   l  L   l  L  �  �  �      F  , ,    �     l  �   l  �  �    �      F  , ,    �     l  �   l  �  �    �      F  , ,  �  �  �   l  l   l  l  �  �  �      F  , ,  �  �  �   l  l   l  l  �  �  �      F  , ,  	�  !4  	�  !�  
�  !�  
�  !4  	�  !4      F  , ,  	�  !4  	�  !�  
�  !�  
�  !4  	�  !4      F  , ,  �  "�  �  #�  l  #�  l  "�  �  "�      F  , ,  �  "�  �  #�  l  #�  l  "�  �  "�      F  , ,  �  !4  �  !�  L  !�  L  !4  �  !4      F  , ,  �  !4  �  !�  L  !�  L  !4  �  !4      F  , ,  �  $T  �  %  L  %  L  $T  �  $T      F  , ,  �  $T  �  %  L  %  L  $T  �  $T      F  , ,    $T    %  �  %  �  $T    $T      F  , ,    $T    %  �  %  �  $T    $T      F  , ,  �  $T  �  %  l  %  l  $T  �  $T      F  , ,  �  $T  �  %  l  %  l  $T  �  $T      F  , ,  4  �  4   l  �   l  �  �  4  �      F  , ,  4  �  4   l  �   l  �  �  4  �      F  , ,  	�  �  	�   l  
�   l  
�  �  	�  �      F  , ,  	�  �  	�   l  
�   l  
�  �  	�  �      F  , ,  �  %�  �  &�  L  &�  L  %�  �  %�      F  , ,  �  %�  �  &�  L  &�  L  %�  �  %�      F  , ,    %�    &�  �  &�  �  %�    %�      F  , ,    %�    &�  �  &�  �  %�    %�      F  , ,  �  %�  �  &�  l  &�  l  %�  �  %�      F  , ,  �  %�  �  &�  l  &�  l  %�  �  %�      F  , ,  4  %�  4  &�  �  &�  �  %�  4  %�      F  , ,  4  %�  4  &�  �  &�  �  %�  4  %�      F  , ,  	�  %�  	�  &�  
�  &�  
�  %�  	�  %�      F  , ,  	�  %�  	�  &�  
�  &�  
�  %�  	�  %�      F  , ,  	�  "�  	�  #�  
�  #�  
�  "�  	�  "�      F  , ,  	�  "�  	�  #�  
�  #�  
�  "�  	�  "�      F  , ,  T  !4  T  !�    !�    !4  T  !4      F  , ,  T  !4  T  !�    !�    !4  T  !4      F  , ,  �  !4  �  !�  �  !�  �  !4  �  !4      F  , ,  �  !4  �  !�  �  !�  �  !4  �  !4      F  , ,  T  $T  T  %    %    $T  T  $T      F  , ,  T  $T  T  %    %    $T  T  $T      F  , ,  �  $T  �  %  �  %  �  $T  �  $T      F  , ,  �  $T  �  %  �  %  �  $T  �  $T      F  , ,  t  $T  t  %  <  %  <  $T  t  $T      F  , ,  t  $T  t  %  <  %  <  $T  t  $T      F  , ,    $T    %  �  %  �  $T    $T      F  , ,    $T    %  �  %  �  $T    $T      F  , ,  �  $T  �  %  \  %  \  $T  �  $T      F  , ,  �  $T  �  %  \  %  \  $T  �  $T      F  , ,  t  !4  t  !�  <  !�  <  !4  t  !4      F  , ,  t  !4  t  !�  <  !�  <  !4  t  !4      F  , ,    !4    !�  �  !�  �  !4    !4      F  , ,    !4    !�  �  !�  �  !4    !4      F  , ,  T  �  T   l     l    �  T  �      F  , ,  T  �  T   l     l    �  T  �      F  , ,  �  �  �   l  �   l  �  �  �  �      F  , ,  �  �  �   l  �   l  �  �  �  �      F  , ,  t  �  t   l  <   l  <  �  t  �      F  , ,  t  �  t   l  <   l  <  �  t  �      F  , ,    �     l  �   l  �  �    �      F  , ,    �     l  �   l  �  �    �      F  , ,  �  �  �   l  \   l  \  �  �  �      F  , ,  �  �  �   l  \   l  \  �  �  �      F  , ,  t  "�  t  #�  <  #�  <  "�  t  "�      F  , ,  t  "�  t  #�  <  #�  <  "�  t  "�      F  , ,    "�    #�  �  #�  �  "�    "�      F  , ,    "�    #�  �  #�  �  "�    "�      F  , ,  �  %�  �  &�  \  &�  \  %�  �  %�      F  , ,  �  %�  �  &�  \  &�  \  %�  �  %�      F  , ,  �  !4  �  !�  \  !�  \  !4  �  !4      F  , ,  �  !4  �  !�  \  !�  \  !4  �  !4      F  , ,  �  "�  �  #�  \  #�  \  "�  �  "�      F  , ,  �  "�  �  #�  \  #�  \  "�  �  "�      F  , ,  T  %�  T  &�    &�    %�  T  %�      F  , ,  T  %�  T  &�    &�    %�  T  %�      F  , ,  �  %�  �  &�  �  &�  �  %�  �  %�      F  , ,  �  %�  �  &�  �  &�  �  %�  �  %�      F  , ,  t  %�  t  &�  <  &�  <  %�  t  %�      F  , ,  t  %�  t  &�  <  &�  <  %�  t  %�      F  , ,    %�    &�  �  &�  �  %�    %�      F  , ,    %�    &�  �  &�  �  %�    %�      F  , ,  �  "�  �  #�  �  #�  �  "�  �  "�      F  , ,  �  "�  �  #�  �  #�  �  "�  �  "�      F  , ,  T  "�  T  #�    #�    "�  T  "�      F  , ,  T  "�  T  #�    #�    "�  T  "�      F  , ,  d  't  d  (<  ,  (<  ,  't  d  't      F  , ,  d  't  d  (<  ,  (<  ,  't  d  't      F  , ,  d  $T  d  %  ,  %  ,  $T  d  $T      F  , ,  d  $T  d  %  ,  %  ,  $T  d  $T      F  , ,  d  )  d  )�  ,  )�  ,  )  d  )      F  , ,  d  )  d  )�  ,  )�  ,  )  d  )      F  , ,  d  "�  d  #�  ,  #�  ,  "�  d  "�      F  , ,  d  "�  d  #�  ,  #�  ,  "�  d  "�      F  , ,  d  %�  d  &�  ,  &�  ,  %�  d  %�      F  , ,  d  %�  d  &�  ,  &�  ,  %�  d  %�      F  , ,  d  ,$  d  ,�  ,  ,�  ,  ,$  d  ,$      F  , ,  d  ,$  d  ,�  ,  ,�  ,  ,$  d  ,$      F  , ,  d  *�  d  +\  ,  +\  ,  *�  d  *�      F  , ,  d  *�  d  +\  ,  +\  ,  *�  d  *�      F  , ,  d  �  d   l  ,   l  ,  �  d  �      F  , ,  d  �  d   l  ,   l  ,  �  d  �      F  , ,  d  !4  d  !�  ,  !�  ,  !4  d  !4      F  , ,  d  !4  d  !�  ,  !�  ,  !4  d  !4      F  , ,  �  )  �  )�   l  )�   l  )  �  )      F  , ,  �  )  �  )�   l  )�   l  )  �  )      F  , ,  �  't  �  (<   l  (<   l  't  �  't      F  , ,  �  't  �  (<   l  (<   l  't  �  't      F  , ,  �  't  �  (<  L  (<  L  't  �  't      F  , ,  �  't  �  (<  L  (<  L  't  �  't      F  , ,    't    (<  �  (<  �  't    't      F  , ,    't    (<  �  (<  �  't    't      F  , ,  �  't  �  (<  �  (<  �  't  �  't      F  , ,  �  't  �  (<  �  (<  �  't  �  't      F  , ,  �  ,$  �  ,�  �  ,�  �  ,$  �  ,$      F  , ,  �  ,$  �  ,�  �  ,�  �  ,$  �  ,$      F  , ,  �  ,$  �  ,�  L  ,�  L  ,$  �  ,$      F  , ,  �  ,$  �  ,�  L  ,�  L  ,$  �  ,$      F  , ,    ,$    ,�  �  ,�  �  ,$    ,$      F  , ,    ,$    ,�  �  ,�  �  ,$    ,$      F  , ,  �  ,$  �  ,�   l  ,�   l  ,$  �  ,$      F  , ,  �  ,$  �  ,�   l  ,�   l  ,$  �  ,$      F  , ,  �  )  �  )�  �  )�  �  )  �  )      F  , ,  �  )  �  )�  �  )�  �  )  �  )      F  , ,  �  *�  �  +\  �  +\  �  *�  �  *�      F  , ,  �  *�  �  +\  �  +\  �  *�  �  *�      F  , ,  �  *�  �  +\  L  +\  L  *�  �  *�      F  , ,  �  *�  �  +\  L  +\  L  *�  �  *�      F  , ,    *�    +\  �  +\  �  *�    *�      F  , ,    *�    +\  �  +\  �  *�    *�      F  , ,  �  *�  �  +\   l  +\   l  *�  �  *�      F  , ,  �  *�  �  +\   l  +\   l  *�  �  *�      F  , ,  �  )  �  )�  L  )�  L  )  �  )      F  , ,  �  )  �  )�  L  )�  L  )  �  )      F  , ,    )    )�  �  )�  �  )    )      F  , ,    )    )�  �  )�  �  )    )      F  , ,  D  ,$  D  ,�    ,�    ,$  D  ,$      F  , ,  D  ,$  D  ,�    ,�    ,$  D  ,$      F  , ,  �  ,$  �  ,�  �  ,�  �  ,$  �  ,$      F  , ,  �  ,$  �  ,�  �  ,�  �  ,$  �  ,$      F  , ,  �  't  �  (<  |  (<  |  't  �  't      F  , ,  �  't  �  (<  |  (<  |  't  �  't      F  , ,  D  't  D  (<    (<    't  D  't      F  , ,  D  't  D  (<    (<    't  D  't      F  , ,  $  )  $  )�  �  )�  �  )  $  )      F  , ,  $  )  $  )�  �  )�  �  )  $  )      F  , ,  �  )  �  )�  |  )�  |  )  �  )      F  , ,  �  )  �  )�  |  )�  |  )  �  )      F  , ,  D  )  D  )�    )�    )  D  )      F  , ,  D  )  D  )�    )�    )  D  )      F  , ,  �  *�  �  +\  �  +\  �  *�  �  *�      F  , ,  �  *�  �  +\  �  +\  �  *�  �  *�      F  , ,  �  )  �  )�  �  )�  �  )  �  )      F  , ,  �  )  �  )�  �  )�  �  )  �  )      F  , ,  �  't  �  (<  �  (<  �  't  �  't      F  , ,  �  't  �  (<  �  (<  �  't  �  't      F  , ,  $  *�  $  +\  �  +\  �  *�  $  *�      F  , ,  $  *�  $  +\  �  +\  �  *�  $  *�      F  , ,  �  *�  �  +\  |  +\  |  *�  �  *�      F  , ,  �  *�  �  +\  |  +\  |  *�  �  *�      F  , ,  D  *�  D  +\    +\    *�  D  *�      F  , ,  D  *�  D  +\    +\    *�  D  *�      F  , ,  $  ,$  $  ,�  �  ,�  �  ,$  $  ,$      F  , ,  $  ,$  $  ,�  �  ,�  �  ,$  $  ,$      F  , ,  �  ,$  �  ,�  |  ,�  |  ,$  �  ,$      F  , ,  �  ,$  �  ,�  |  ,�  |  ,$  �  ,$      F  , ,  $  't  $  (<  �  (<  �  't  $  't      F  , ,  $  't  $  (<  �  (<  �  't  $  't      F  , ,  $  !4  $  !�  �  !�  �  !4  $  !4      F  , ,  $  !4  $  !�  �  !�  �  !4  $  !4      F  , ,  �  !4  �  !�  |  !�  |  !4  �  !4      F  , ,  �  !4  �  !�  |  !�  |  !4  �  !4      F  , ,  �  "�  �  #�  �  #�  �  "�  �  "�      F  , ,  �  "�  �  #�  �  #�  �  "�  �  "�      F  , ,  �  $T  �  %  �  %  �  $T  �  $T      F  , ,  �  $T  �  %  �  %  �  $T  �  $T      F  , ,  $  "�  $  #�  �  #�  �  "�  $  "�      F  , ,  $  "�  $  #�  �  #�  �  "�  $  "�      F  , ,  �  "�  �  #�  |  #�  |  "�  �  "�      F  , ,  �  "�  �  #�  |  #�  |  "�  �  "�      F  , ,  D  "�  D  #�    #�    "�  D  "�      F  , ,  D  "�  D  #�    #�    "�  D  "�      F  , ,  �  $T  �  %  |  %  |  $T  �  $T      F  , ,  �  $T  �  %  |  %  |  $T  �  $T      F  , ,  $  �  $   l  �   l  �  �  $  �      F  , ,  $  �  $   l  �   l  �  �  $  �      F  , ,  �  �  �   l  |   l  |  �  �  �      F  , ,  �  �  �   l  |   l  |  �  �  �      F  , ,  D  �  D   l     l    �  D  �      F  , ,  D  �  D   l     l    �  D  �      F  , ,  �  �  �   l  �   l  �  �  �  �      F  , ,  �  �  �   l  �   l  �  �  �  �      F  , ,  �  %�  �  &�  �  &�  �  %�  �  %�      F  , ,  �  %�  �  &�  �  &�  �  %�  �  %�      F  , ,  $  %�  $  &�  �  &�  �  %�  $  %�      F  , ,  $  %�  $  &�  �  &�  �  %�  $  %�      F  , ,  D  !4  D  !�    !�    !4  D  !4      F  , ,  D  !4  D  !�    !�    !4  D  !4      F  , ,  �  !4  �  !�  �  !�  �  !4  �  !4      F  , ,  �  !4  �  !�  �  !�  �  !4  �  !4      F  , ,  $  $T  $  %  �  %  �  $T  $  $T      F  , ,  $  $T  $  %  �  %  �  $T  $  $T      F  , ,  �  %�  �  &�  |  &�  |  %�  �  %�      F  , ,  �  %�  �  &�  |  &�  |  %�  �  %�      F  , ,  D  %�  D  &�    &�    %�  D  %�      F  , ,  D  %�  D  &�    &�    %�  D  %�      F  , ,  D  $T  D  %    %    $T  D  $T      F  , ,  D  $T  D  %    %    $T  D  $T      F  , ,  �  $T  �  %  L  %  L  $T  �  $T      F  , ,  �  $T  �  %  L  %  L  $T  �  $T      F  , ,    $T    %  �  %  �  $T    $T      F  , ,    $T    %  �  %  �  $T    $T      F  , ,  �  $T  �  %   l  %   l  $T  �  $T      F  , ,  �  $T  �  %   l  %   l  $T  �  $T      F  , ,  �  !4  �  !�  �  !�  �  !4  �  !4      F  , ,  �  !4  �  !�  �  !�  �  !4  �  !4      F  , ,  �  !4  �  !�  L  !�  L  !4  �  !4      F  , ,  �  !4  �  !�  L  !�  L  !4  �  !4      F  , ,  �  %�  �  &�  �  &�  �  %�  �  %�      F  , ,  �  %�  �  &�  �  &�  �  %�  �  %�      F  , ,  �  %�  �  &�  L  &�  L  %�  �  %�      F  , ,  �  %�  �  &�  L  &�  L  %�  �  %�      F  , ,    %�    &�  �  &�  �  %�    %�      F  , ,    %�    &�  �  &�  �  %�    %�      F  , ,  �  %�  �  &�   l  &�   l  %�  �  %�      F  , ,  �  %�  �  &�   l  &�   l  %�  �  %�      F  , ,    !4    !�  �  !�  �  !4    !4      F  , ,    !4    !�  �  !�  �  !4    !4      F  , ,  �  !4  �  !�   l  !�   l  !4  �  !4      F  , ,  �  !4  �  !�   l  !�   l  !4  �  !4      F  , ,    �     l  �   l  �  �    �      F  , ,    �     l  �   l  �  �    �      F  , ,  �  �  �   l   l   l   l  �  �  �      F  , ,  �  �  �   l   l   l   l  �  �  �      F  , ,  �  "�  �  #�   l  #�   l  "�  �  "�      F  , ,  �  "�  �  #�   l  #�   l  "�  �  "�      F  , ,  �  �  �   l  �   l  �  �  �  �      F  , ,  �  �  �   l  �   l  �  �  �  �      F  , ,  �  �  �   l  L   l  L  �  �  �      F  , ,  �  �  �   l  L   l  L  �  �  �      F  , ,  �  $T  �  %  �  %  �  $T  �  $T      F  , ,  �  $T  �  %  �  %  �  $T  �  $T      F  , ,  �  "�  �  #�  �  #�  �  "�  �  "�      F  , ,  �  "�  �  #�  �  #�  �  "�  �  "�      F  , ,  �  "�  �  #�  L  #�  L  "�  �  "�      F  , ,  �  "�  �  #�  L  #�  L  "�  �  "�      F  , ,    "�    #�  �  #�  �  "�    "�      F  , ,    "�    #�  �  #�  �  "�    "�      F  , ,  �    �  �  L  �  L    �        F  , ,  �    �  �  L  �  L    �        F  , ,        �  �  �  �            F  , ,        �  �  �  �            F  , ,  �    �  �  l  �  l    �        F  , ,  �    �  �  l  �  l    �        F  , ,  4    4  �  �  �  �    4        F  , ,  4    4  �  �  �  �    4        F  , ,  	�    	�  �  
�  �  
�    	�        F  , ,  	�    	�  �  
�  �  
�    	�        F  , ,  T    T  �    �      T        F  , ,  T    T  �    �      T        F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  �  �  �    �        F  , ,  t    t  �  <  �  <    t        F  , ,  t    t  �  <  �  <    t        F  , ,        �  �  �  �            F  , ,        �  �  �  �            F  , ,  �    �  �  \  �  \    �        F  , ,  �    �  �  \  �  \    �        F  , ,  $    $  �  �  �  �    $        F  , ,  $    $  �  �  �  �    $        F  , ,  �    �  �  |  �  |    �        F  , ,  �    �  �  |  �  |    �        F  , ,  D    D  �    �      D        F  , ,  D    D  �    �      D        F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  �  �  �    �        F  , ,  d    d  �  ,  �  ,    d        F  , ,  d    d  �  ,  �  ,    d        F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  L  �  L    �        F  , ,  �    �  �  L  �  L    �        F  , ,        �  �  �  �            F  , ,        �  �  �  �            F  , ,  �    �  �   l  �   l    �        F  , ,  �    �  �   l  �   l    �        F  , ,  d    d  �  ,  �  ,    d        F  , ,  d    d  �  ,  �  ,    d        F  , ,  d  �  d  \  ,  \  ,  �  d  �      F  , ,  d  �  d  \  ,  \  ,  �  d  �      F  , ,  d  $  d  �  ,  �  ,  $  d  $      F  , ,  d  $  d  �  ,  �  ,  $  d  $      F  , ,  d  �  d  |  ,  |  ,  �  d  �      F  , ,  d  �  d  |  ,  |  ,  �  d  �      F  , ,  d  D  d    ,    ,  D  d  D      F  , ,  d  D  d    ,    ,  D  d  D      F  , ,  d  �  d  �  ,  �  ,  �  d  �      F  , ,  d  �  d  �  ,  �  ,  �  d  �      F  , ,  d  d  d  ,  ,  ,  ,  d  d  d      F  , ,  d  d  d  ,  ,  ,  ,  d  d  d      F  , ,  d  �  d  �  ,  �  ,  �  d  �      F  , ,  d  �  d  �  ,  �  ,  �  d  �      F  , ,  d  �  d  L  ,  L  ,  �  d  �      F  , ,  d  �  d  L  ,  L  ,  �  d  �      F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  �  �  �    �        F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,    �    �  �  �  �  �    �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �   l  �   l  �  �  �      F  , ,  �  �  �  �   l  �   l  �  �  �      F  , ,  �    �  �  L  �  L    �        F  , ,  �    �  �  L  �  L    �        F  , ,  �  d  �  ,  �  ,  �  d  �  d      F  , ,  �  d  �  ,  �  ,  �  d  �  d      F  , ,  �  d  �  ,  L  ,  L  d  �  d      F  , ,  �  d  �  ,  L  ,  L  d  �  d      F  , ,    d    ,  �  ,  �  d    d      F  , ,    d    ,  �  ,  �  d    d      F  , ,  �  d  �  ,   l  ,   l  d  �  d      F  , ,  �  d  �  ,   l  ,   l  d  �  d      F  , ,        �  �  �  �            F  , ,        �  �  �  �            F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,    �    �  �  �  �  �    �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �   l  �   l  �  �  �      F  , ,  �  �  �  �   l  �   l  �  �  �      F  , ,  �    �  �   l  �   l    �        F  , ,  �    �  �   l  �   l    �        F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  �  �  �  L  L  L  L  �  �  �      F  , ,  �  �  �  L  L  L  L  �  �  �      F  , ,    �    L  �  L  �  �    �      F  , ,    �    L  �  L  �  �    �      F  , ,  �  �  �  L   l  L   l  �  �  �      F  , ,  �  �  �  L   l  L   l  �  �  �      F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  |  �  |    �        F  , ,  �    �  �  |  �  |    �        F  , ,  $  �  $  �  �  �  �  �  $  �      F  , ,  $  �  $  �  �  �  �  �  $  �      F  , ,  �  �  �  �  |  �  |  �  �  �      F  , ,  �  �  �  �  |  �  |  �  �  �      F  , ,  D  �  D  �    �    �  D  �      F  , ,  D  �  D  �    �    �  D  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  D    D  �    �      D        F  , ,  D    D  �    �      D        F  , ,  $    $  �  �  �  �    $        F  , ,  $    $  �  �  �  �    $        F  , ,  $  �  $  �  �  �  �  �  $  �      F  , ,  $  �  $  �  �  �  �  �  $  �      F  , ,  $  d  $  ,  �  ,  �  d  $  d      F  , ,  $  d  $  ,  �  ,  �  d  $  d      F  , ,  �  d  �  ,  |  ,  |  d  �  d      F  , ,  �  d  �  ,  |  ,  |  d  �  d      F  , ,  $  �  $  L  �  L  �  �  $  �      F  , ,  $  �  $  L  �  L  �  �  $  �      F  , ,  �  �  �  L  |  L  |  �  �  �      F  , ,  �  �  �  L  |  L  |  �  �  �      F  , ,  D  �  D  L    L    �  D  �      F  , ,  D  �  D  L    L    �  D  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  D  d  D  ,    ,    d  D  d      F  , ,  D  d  D  ,    ,    d  D  d      F  , ,  �  d  �  ,  �  ,  �  d  �  d      F  , ,  �  d  �  ,  �  ,  �  d  �  d      F  , ,  �  �  �  �  |  �  |  �  �  �      F  , ,  �  �  �  �  |  �  |  �  �  �      F  , ,  D  �  D  �    �    �  D  �      F  , ,  D  �  D  �    �    �  D  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  $  �  �  �  �  �  $  �  $      F  , ,  �  $  �  �  �  �  �  $  �  $      F  , ,  �  �  �  \  |  \  |  �  �  �      F  , ,  �  �  �  \  |  \  |  �  �  �      F  , ,  $  �  $  |  �  |  �  �  $  �      F  , ,  $  �  $  |  �  |  �  �  $  �      F  , ,  �  �  �  |  |  |  |  �  �  �      F  , ,  �  �  �  |  |  |  |  �  �  �      F  , ,  D  �  D  |    |    �  D  �      F  , ,  D  �  D  |    |    �  D  �      F  , ,  �  �  �  |  �  |  �  �  �  �      F  , ,  �  �  �  |  �  |  �  �  �  �      F  , ,  D  �  D  \    \    �  D  �      F  , ,  D  �  D  \    \    �  D  �      F  , ,  $  D  $    �    �  D  $  D      F  , ,  $  D  $    �    �  D  $  D      F  , ,  �  D  �    |    |  D  �  D      F  , ,  �  D  �    |    |  D  �  D      F  , ,  D  D  D          D  D  D      F  , ,  D  D  D          D  D  D      F  , ,  �  D  �    �    �  D  �  D      F  , ,  �  D  �    �    �  D  �  D      F  , ,  �  �  �  \  �  \  �  �  �  �      F  , ,  �  �  �  \  �  \  �  �  �  �      F  , ,  $  �  $  \  �  \  �  �  $  �      F  , ,  $  �  $  \  �  \  �  �  $  �      F  , ,  $  $  $  �  �  �  �  $  $  $      F  , ,  $  $  $  �  �  �  �  $  $  $      F  , ,  �  $  �  �  |  �  |  $  �  $      F  , ,  �  $  �  �  |  �  |  $  �  $      F  , ,  D  $  D  �    �    $  D  $      F  , ,  D  $  D  �    �    $  D  $      F  , ,  �  �  �  |  L  |  L  �  �  �      F  , ,  �  �  �  |  L  |  L  �  �  �      F  , ,    �    |  �  |  �  �    �      F  , ,    �    |  �  |  �  �    �      F  , ,  �  �  �  |   l  |   l  �  �  �      F  , ,  �  �  �  |   l  |   l  �  �  �      F  , ,  �  $  �  �  L  �  L  $  �  $      F  , ,  �  $  �  �  L  �  L  $  �  $      F  , ,    $    �  �  �  �  $    $      F  , ,    $    �  �  �  �  $    $      F  , ,  �  $  �  �   l  �   l  $  �  $      F  , ,  �  $  �  �   l  �   l  $  �  $      F  , ,  �  �  �  \  L  \  L  �  �  �      F  , ,  �  �  �  \  L  \  L  �  �  �      F  , ,    �    \  �  \  �  �    �      F  , ,    �    \  �  \  �  �    �      F  , ,  �  D  �    �    �  D  �  D      F  , ,  �  D  �    �    �  D  �  D      F  , ,  �  D  �    L    L  D  �  D      F  , ,  �  D  �    L    L  D  �  D      F  , ,    D      �    �  D    D      F  , ,    D      �    �  D    D      F  , ,  �  D  �     l     l  D  �  D      F  , ,  �  D  �     l     l  D  �  D      F  , ,  �  �  �  \   l  \   l  �  �  �      F  , ,  �  �  �  \   l  \   l  �  �  �      F  , ,  �  �  �  \  �  \  �  �  �  �      F  , ,  �  �  �  \  �  \  �  �  �  �      F  , ,  �  $  �  �  �  �  �  $  �  $      F  , ,  �  $  �  �  �  �  �  $  �  $      F  , ,  �  �  �  |  �  |  �  �  �  �      F  , ,  �  �  �  |  �  |  �  �  �  �      F  , ,  T  �  T  �    �    �  T  �      F  , ,  T  �  T  �    �    �  T  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  t  �  t  �  <  �  <  �  t  �      F  , ,  t  �  t  �  <  �  <  �  t  �      F  , ,    �    �  �  �  �  �    �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  \  �  \  �  �  �      F  , ,  �  �  �  �  \  �  \  �  �  �      F  , ,        �  �  �  �            F  , ,        �  �  �  �            F  , ,  �    �  �  \  �  \    �        F  , ,  �    �  �  \  �  \    �        F  , ,  T  d  T  ,    ,    d  T  d      F  , ,  T  d  T  ,    ,    d  T  d      F  , ,  �  d  �  ,  �  ,  �  d  �  d      F  , ,  �  d  �  ,  �  ,  �  d  �  d      F  , ,  t  d  t  ,  <  ,  <  d  t  d      F  , ,  t  d  t  ,  <  ,  <  d  t  d      F  , ,    d    ,  �  ,  �  d    d      F  , ,    d    ,  �  ,  �  d    d      F  , ,  �  d  �  ,  \  ,  \  d  �  d      F  , ,  �  d  �  ,  \  ,  \  d  �  d      F  , ,  T  �  T  �    �    �  T  �      F  , ,  T  �  T  �    �    �  T  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  t  �  t  �  <  �  <  �  t  �      F  , ,  t  �  t  �  <  �  <  �  t  �      F  , ,    �    �  �  �  �  �    �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  \  �  \  �  �  �      F  , ,  �  �  �  �  \  �  \  �  �  �      F  , ,  T    T  �    �      T        F  , ,  T    T  �    �      T        F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  �  �  �    �        F  , ,  t    t  �  <  �  <    t        F  , ,  t    t  �  <  �  <    t        F  , ,  T  �  T  L    L    �  T  �      F  , ,  T  �  T  L    L    �  T  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  t  �  t  L  <  L  <  �  t  �      F  , ,  t  �  t  L  <  L  <  �  t  �      F  , ,    �    L  �  L  �  �    �      F  , ,    �    L  �  L  �  �    �      F  , ,  �  �  �  L  \  L  \  �  �  �      F  , ,  �  �  �  L  \  L  \  �  �  �      F  , ,  4  �  4  �  �  �  �  �  4  �      F  , ,  4  �  4  �  �  �  �  �  4  �      F  , ,  	�  �  	�  �  
�  �  
�  �  	�  �      F  , ,  	�  �  	�  �  
�  �  
�  �  	�  �      F  , ,  �  d  �  ,  L  ,  L  d  �  d      F  , ,  �  d  �  ,  L  ,  L  d  �  d      F  , ,    d    ,  �  ,  �  d    d      F  , ,    d    ,  �  ,  �  d    d      F  , ,  �  d  �  ,  l  ,  l  d  �  d      F  , ,  �  d  �  ,  l  ,  l  d  �  d      F  , ,  4  d  4  ,  �  ,  �  d  4  d      F  , ,  4  d  4  ,  �  ,  �  d  4  d      F  , ,  	�  d  	�  ,  
�  ,  
�  d  	�  d      F  , ,  	�  d  	�  ,  
�  ,  
�  d  	�  d      F  , ,  	�    	�  �  
�  �  
�    	�        F  , ,  	�    	�  �  
�  �  
�    	�        F  , ,  �  �  �  �  l  �  l  �  �  �      F  , ,  �  �  �  �  l  �  l  �  �  �      F  , ,  4  �  4  �  �  �  �  �  4  �      F  , ,  4  �  4  �  �  �  �  �  4  �      F  , ,  	�  �  	�  �  
�  �  
�  �  	�  �      F  , ,  	�  �  	�  �  
�  �  
�  �  	�  �      F  , ,  �  �  �  L  L  L  L  �  �  �      F  , ,  �  �  �  L  L  L  L  �  �  �      F  , ,    �    L  �  L  �  �    �      F  , ,    �    L  �  L  �  �    �      F  , ,  �  �  �  L  l  L  l  �  �  �      F  , ,  �  �  �  L  l  L  l  �  �  �      F  , ,  4  �  4  L  �  L  �  �  4  �      F  , ,  4  �  4  L  �  L  �  �  4  �      F  , ,  	�  �  	�  L  
�  L  
�  �  	�  �      F  , ,  	�  �  	�  L  
�  L  
�  �  	�  �      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,    �    �  �  �  �  �    �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,    �    �  �  �  �  �    �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  l  �  l  �  �  �      F  , ,  �  �  �  �  l  �  l  �  �  �      F  , ,  �    �  �  L  �  L    �        F  , ,  �    �  �  L  �  L    �        F  , ,        �  �  �  �            F  , ,        �  �  �  �            F  , ,  �    �  �  l  �  l    �        F  , ,  �    �  �  l  �  l    �        F  , ,  4    4  �  �  �  �    4        F  , ,  4    4  �  �  �  �    4        F  , ,    $    �  �  �  �  $    $      F  , ,    $    �  �  �  �  $    $      F  , ,  	�  �  	�  \  
�  \  
�  �  	�  �      F  , ,  	�  �  	�  \  
�  \  
�  �  	�  �      F  , ,  	�  $  	�  �  
�  �  
�  $  	�  $      F  , ,  	�  $  	�  �  
�  �  
�  $  	�  $      F  , ,    �    |  �  |  �  �    �      F  , ,    �    |  �  |  �  �    �      F  , ,  �  �  �  |  l  |  l  �  �  �      F  , ,  �  �  �  |  l  |  l  �  �  �      F  , ,  4  �  4  |  �  |  �  �  4  �      F  , ,  4  �  4  |  �  |  �  �  4  �      F  , ,  	�  �  	�  |  
�  |  
�  �  	�  �      F  , ,  	�  �  	�  |  
�  |  
�  �  	�  �      F  , ,  4  �  4  \  �  \  �  �  4  �      F  , ,  4  �  4  \  �  \  �  �  4  �      F  , ,  �  �  �  |  L  |  L  �  �  �      F  , ,  �  �  �  |  L  |  L  �  �  �      F  , ,  �  $  �  �  l  �  l  $  �  $      F  , ,  �  $  �  �  l  �  l  $  �  $      F  , ,  4  $  4  �  �  �  �  $  4  $      F  , ,  4  $  4  �  �  �  �  $  4  $      F  , ,  �  D  �    L    L  D  �  D      F  , ,  �  D  �    L    L  D  �  D      F  , ,    D      �    �  D    D      F  , ,    D      �    �  D    D      F  , ,  �  D  �    l    l  D  �  D      F  , ,  �  D  �    l    l  D  �  D      F  , ,  4  D  4    �    �  D  4  D      F  , ,  4  D  4    �    �  D  4  D      F  , ,  	�  D  	�    
�    
�  D  	�  D      F  , ,  	�  D  	�    
�    
�  D  	�  D      F  , ,  �  �  �  \  L  \  L  �  �  �      F  , ,  �  �  �  \  L  \  L  �  �  �      F  , ,    �    \  �  \  �  �    �      F  , ,    �    \  �  \  �  �    �      F  , ,  �  �  �  \  l  \  l  �  �  �      F  , ,  �  �  �  \  l  \  l  �  �  �      F  , ,  �  $  �  �  L  �  L  $  �  $      F  , ,  �  $  �  �  L  �  L  $  �  $      F  , ,  T  $  T  �    �    $  T  $      F  , ,  T  $  T  �    �    $  T  $      F  , ,  �  $  �  �  �  �  �  $  �  $      F  , ,  �  $  �  �  �  �  �  $  �  $      F  , ,  t  $  t  �  <  �  <  $  t  $      F  , ,  t  $  t  �  <  �  <  $  t  $      F  , ,    $    �  �  �  �  $    $      F  , ,    $    �  �  �  �  $    $      F  , ,  �  $  �  �  \  �  \  $  �  $      F  , ,  �  $  �  �  \  �  \  $  �  $      F  , ,  T  �  T  |    |    �  T  �      F  , ,  T  �  T  |    |    �  T  �      F  , ,  �  �  �  |  �  |  �  �  �  �      F  , ,  �  �  �  |  �  |  �  �  �  �      F  , ,  t  �  t  |  <  |  <  �  t  �      F  , ,  t  �  t  |  <  |  <  �  t  �      F  , ,    �    |  �  |  �  �    �      F  , ,    �    |  �  |  �  �    �      F  , ,  �  �  �  |  \  |  \  �  �  �      F  , ,  �  �  �  |  \  |  \  �  �  �      F  , ,  T  �  T  \    \    �  T  �      F  , ,  T  �  T  \    \    �  T  �      F  , ,  �  �  �  \  �  \  �  �  �  �      F  , ,  �  �  �  \  �  \  �  �  �  �      F  , ,  T  D  T          D  T  D      F  , ,  T  D  T          D  T  D      F  , ,  �  D  �    �    �  D  �  D      F  , ,  �  D  �    �    �  D  �  D      F  , ,  t  D  t    <    <  D  t  D      F  , ,  t  D  t    <    <  D  t  D      F  , ,    D      �    �  D    D      F  , ,    D      �    �  D    D      F  , ,  t  �  t  \  <  \  <  �  t  �      F  , ,  t  �  t  \  <  \  <  �  t  �      F  , ,    �    \  �  \  �  �    �      F  , ,    �    \  �  \  �  �    �      F  , ,  �  �  �  \  \  \  \  �  �  �      F  , ,  �  �  �  \  \  \  \  �  �  �      F  , ,  �  D  �    \    \  D  �  D      F  , ,  �  D  �    \    \  D  �  D      F  , ,  �  4  �  �  L  �  L  4  �  4      F  , ,  �  4  �  �  L  �  L  4  �  4      F  , ,    4    �  �  �  �  4    4      F  , ,    4    �  �  �  �  4    4      F  , ,  �  4  �  �  l  �  l  4  �  4      F  , ,  �  4  �  �  l  �  l  4  �  4      F  , ,  4  4  4  �  �  �  �  4  4  4      F  , ,  4  4  4  �  �  �  �  4  4  4      F  , ,  	�  4  	�  �  
�  �  
�  4  	�  4      F  , ,  	�  4  	�  �  
�  �  
�  4  	�  4      F  , ,  T  4  T  �    �    4  T  4      F  , ,  T  4  T  �    �    4  T  4      F  , ,  �  4  �  �  �  �  �  4  �  4      F  , ,  �  4  �  �  �  �  �  4  �  4      F  , ,  t  4  t  �  <  �  <  4  t  4      F  , ,  t  4  t  �  <  �  <  4  t  4      F  , ,    4    �  �  �  �  4    4      F  , ,    4    �  �  �  �  4    4      F  , ,  �  4  �  �  \  �  \  4  �  4      F  , ,  �  4  �  �  \  �  \  4  �  4      F  , ,  T  	�  T  
�    
�    	�  T  	�      F  , ,  T  	�  T  
�    
�    	�  T  	�      F  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      F  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      F  , ,  t  	�  t  
�  <  
�  <  	�  t  	�      F  , ,  t  	�  t  
�  <  
�  <  	�  t  	�      F  , ,    	�    
�  �  
�  �  	�    	�      F  , ,    	�    
�  �  
�  �  	�    	�      F  , ,  �  	�  �  
�  \  
�  \  	�  �  	�      F  , ,  �  	�  �  
�  \  
�  \  	�  �  	�      F  , ,  T  T  T          T  T  T      F  , ,  T  T  T          T  T  T      F  , ,  �  T  �    �    �  T  �  T      F  , ,  �  T  �    �    �  T  �  T      F  , ,  t  T  t    <    <  T  t  T      F  , ,  t  T  t    <    <  T  t  T      F  , ,    T      �    �  T    T      F  , ,    T      �    �  T    T      F  , ,  �  T  �    \    \  T  �  T      F  , ,  �  T  �    \    \  T  �  T      F  , ,  T  �  T  �    �    �  T  �      F  , ,  T  �  T  �    �    �  T  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  t  �  t  �  <  �  <  �  t  �      F  , ,  t  �  t  �  <  �  <  �  t  �      F  , ,    �    �  �  �  �  �    �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  \  �  \  �  �  �      F  , ,  �  �  �  �  \  �  \  �  �  �      F  , ,  T  t  T  <    <    t  T  t      F  , ,  T  t  T  <    <    t  T  t      F  , ,  �  t  �  <  �  <  �  t  �  t      F  , ,  �  t  �  <  �  <  �  t  �  t      F  , ,  t  t  t  <  <  <  <  t  t  t      F  , ,  t  t  t  <  <  <  <  t  t  t      F  , ,    t    <  �  <  �  t    t      F  , ,    t    <  �  <  �  t    t      F  , ,  �  t  �  <  \  <  \  t  �  t      F  , ,  �  t  �  <  \  <  \  t  �  t      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,    �    �  �  �  �  �    �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  l  �  l  �  �  �      F  , ,  �  �  �  �  l  �  l  �  �  �      F  , ,  4  �  4  �  �  �  �  �  4  �      F  , ,  4  �  4  �  �  �  �  �  4  �      F  , ,  	�  �  	�  �  
�  �  
�  �  	�  �      F  , ,  	�  �  	�  �  
�  �  
�  �  	�  �      F  , ,  �  T  �    L    L  T  �  T      F  , ,  �  T  �    L    L  T  �  T      F  , ,    T      �    �  T    T      F  , ,    T      �    �  T    T      F  , ,  �  T  �    l    l  T  �  T      F  , ,  �  T  �    l    l  T  �  T      F  , ,  4  T  4    �    �  T  4  T      F  , ,  4  T  4    �    �  T  4  T      F  , ,  	�  T  	�    
�    
�  T  	�  T      F  , ,  	�  T  	�    
�    
�  T  	�  T      F  , ,  �  t  �  <  L  <  L  t  �  t      F  , ,  �  t  �  <  L  <  L  t  �  t      F  , ,    t    <  �  <  �  t    t      F  , ,    t    <  �  <  �  t    t      F  , ,  �  t  �  <  l  <  l  t  �  t      F  , ,  �  t  �  <  l  <  l  t  �  t      F  , ,  4  t  4  <  �  <  �  t  4  t      F  , ,  4  t  4  <  �  <  �  t  4  t      F  , ,  	�  t  	�  <  
�  <  
�  t  	�  t      F  , ,  	�  t  	�  <  
�  <  
�  t  	�  t      F  , ,  �  	�  �  
�  L  
�  L  	�  �  	�      F  , ,  �  	�  �  
�  L  
�  L  	�  �  	�      F  , ,    	�    
�  �  
�  �  	�    	�      F  , ,    	�    
�  �  
�  �  	�    	�      F  , ,  �  	�  �  
�  l  
�  l  	�  �  	�      F  , ,  �  	�  �  
�  l  
�  l  	�  �  	�      F  , ,  4  	�  4  
�  �  
�  �  	�  4  	�      F  , ,  4  	�  4  
�  �  
�  �  	�  4  	�      F  , ,  	�  	�  	�  
�  
�  
�  
�  	�  	�  	�      F  , ,  	�  	�  	�  
�  
�  
�  
�  	�  	�  	�      F  , ,  �  �  �  L  l  L  l  �  �  �      F  , ,  �  �  �  L  l  L  l  �  �  �      F  , ,  4  �  4  L  �  L  �  �  4  �      F  , ,  4  �  4  L  �  L  �  �  4  �      F  , ,  	�  �  	�  L  
�  L  
�  �  	�  �      F  , ,  	�  �  	�  L  
�  L  
�  �  	�  �      F  , ,  �  �  �  L  L  L  L  �  �  �      F  , ,  �  �  �  L  L  L  L  �  �  �      F  , ,  �    �  �  L  �  L    �        F  , ,  �    �  �  L  �  L    �        F  , ,        �  �  �  �            F  , ,        �  �  �  �            F  , ,  �    �  �  l  �  l    �        F  , ,  �    �  �  l  �  l    �        F  , ,  4    4  �  �  �  �    4        F  , ,  4    4  �  �  �  �    4        F  , ,  	�    	�  �  
�  �  
�    	�        F  , ,  	�    	�  �  
�  �  
�    	�        F  , ,    �    L  �  L  �  �    �      F  , ,    �    L  �  L  �  �    �      F  , ,  �  �  �  l  L  l  L  �  �  �      F  , ,  �  �  �  l  L  l  L  �  �  �      F  , ,    �    l  �  l  �  �    �      F  , ,    �    l  �  l  �  �    �      F  , ,  �  �  �  l  l  l  l  �  �  �      F  , ,  �  �  �  l  l  l  l  �  �  �      F  , ,  4  �  4  l  �  l  �  �  4  �      F  , ,  4  �  4  l  �  l  �  �  4  �      F  , ,  	�  �  	�  l  
�  l  
�  �  	�  �      F  , ,  	�  �  	�  l  
�  l  
�  �  	�  �      F  , ,  �  �  �  l  \  l  \  �  �  �      F  , ,  �  �  �  l  \  l  \  �  �  �      F  , ,  T  �  T  l    l    �  T  �      F  , ,  T  �  T  l    l    �  T  �      F  , ,  T  �  T  L    L    �  T  �      F  , ,  T  �  T  L    L    �  T  �      F  , ,  �  �  �  l  �  l  �  �  �  �      F  , ,  �  �  �  l  �  l  �  �  �  �      F  , ,  T    T  �    �      T        F  , ,  T    T  �    �      T        F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  �  �  �    �        F  , ,  t    t  �  <  �  <    t        F  , ,  t    t  �  <  �  <    t        F  , ,        �  �  �  �            F  , ,        �  �  �  �            F  , ,  �    �  �  \  �  \    �        F  , ,  �    �  �  \  �  \    �        F  , ,    �    L  �  L  �  �    �      F  , ,    �    L  �  L  �  �    �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  t  �  t  l  <  l  <  �  t  �      F  , ,  t  �  t  l  <  l  <  �  t  �      F  , ,  t  �  t  L  <  L  <  �  t  �      F  , ,  t  �  t  L  <  L  <  �  t  �      F  , ,  �  �  �  L  \  L  \  �  �  �      F  , ,  �  �  �  L  \  L  \  �  �  �      F  , ,    �    l  �  l  �  �    �      F  , ,    �    l  �  l  �  �    �      F  , ,  d  �  d  l  ,  l  ,  �  d  �      F  , ,  d  �  d  l  ,  l  ,  �  d  �      F  , ,  d  t  d  <  ,  <  ,  t  d  t      F  , ,  d  t  d  <  ,  <  ,  t  d  t      F  , ,  d  	�  d  
�  ,  
�  ,  	�  d  	�      F  , ,  d  	�  d  
�  ,  
�  ,  	�  d  	�      F  , ,  d  �  d  L  ,  L  ,  �  d  �      F  , ,  d  �  d  L  ,  L  ,  �  d  �      F  , ,  d    d  �  ,  �  ,    d        F  , ,  d    d  �  ,  �  ,    d        F  , ,  $  4  $  �  �  �  �  4  $  4      F  , ,  $  4  $  �  �  �  �  4  $  4      F  , ,  �  4  �  �  |  �  |  4  �  4      F  , ,  �  4  �  �  |  �  |  4  �  4      F  , ,  d  T  d    ,    ,  T  d  T      F  , ,  d  T  d    ,    ,  T  d  T      F  , ,  D  4  D  �    �    4  D  4      F  , ,  D  4  D  �    �    4  D  4      F  , ,  �  4  �  �  �  �  �  4  �  4      F  , ,  �  4  �  �  �  �  �  4  �  4      F  , ,  d  4  d  �  ,  �  ,  4  d  4      F  , ,  d  4  d  �  ,  �  ,  4  d  4      F  , ,  �  4  �  �  �  �  �  4  �  4      F  , ,  �  4  �  �  �  �  �  4  �  4      F  , ,  �  4  �  �  L  �  L  4  �  4      F  , ,  �  4  �  �  L  �  L  4  �  4      F  , ,    4    �  �  �  �  4    4      F  , ,    4    �  �  �  �  4    4      F  , ,  �  4  �  �   l  �   l  4  �  4      F  , ,  �  4  �  �   l  �   l  4  �  4      F  , ,  d  �  d  �  ,  �  ,  �  d  �      F  , ,  d  �  d  �  ,  �  ,  �  d  �      F  , ,  �  T  �    �    �  T  �  T      F  , ,  �  T  �    �    �  T  �  T      F  , ,  �  T  �    L    L  T  �  T      F  , ,  �  T  �    L    L  T  �  T      F  , ,    T      �    �  T    T      F  , ,    T      �    �  T    T      F  , ,  �  T  �     l     l  T  �  T      F  , ,  �  T  �     l     l  T  �  T      F  , ,  �  	�  �  
�  L  
�  L  	�  �  	�      F  , ,  �  	�  �  
�  L  
�  L  	�  �  	�      F  , ,    	�    
�  �  
�  �  	�    	�      F  , ,    	�    
�  �  
�  �  	�    	�      F  , ,  �  	�  �  
�   l  
�   l  	�  �  	�      F  , ,  �  	�  �  
�   l  
�   l  	�  �  	�      F  , ,  �  t  �  <  L  <  L  t  �  t      F  , ,  �  t  �  <  L  <  L  t  �  t      F  , ,    t    <  �  <  �  t    t      F  , ,    t    <  �  <  �  t    t      F  , ,  �  t  �  <   l  <   l  t  �  t      F  , ,  �  t  �  <   l  <   l  t  �  t      F  , ,  �  t  �  <  �  <  �  t  �  t      F  , ,  �  t  �  <  �  <  �  t  �  t      F  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      F  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,    �    �  �  �  �  �    �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �   l  �   l  �  �  �      F  , ,  �  �  �  �   l  �   l  �  �  �      F  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      F  , ,  �  	�  �  
�  �  
�  �  	�  �  	�      F  , ,  $  t  $  <  �  <  �  t  $  t      F  , ,  $  t  $  <  �  <  �  t  $  t      F  , ,  �  t  �  <  |  <  |  t  �  t      F  , ,  �  t  �  <  |  <  |  t  �  t      F  , ,  $  T  $    �    �  T  $  T      F  , ,  $  T  $    �    �  T  $  T      F  , ,  �  T  �    |    |  T  �  T      F  , ,  �  T  �    |    |  T  �  T      F  , ,  D  T  D          T  D  T      F  , ,  D  T  D          T  D  T      F  , ,  �  T  �    �    �  T  �  T      F  , ,  �  T  �    �    �  T  �  T      F  , ,  $  �  $  �  �  �  �  �  $  �      F  , ,  $  �  $  �  �  �  �  �  $  �      F  , ,  �  �  �  �  |  �  |  �  �  �      F  , ,  �  �  �  �  |  �  |  �  �  �      F  , ,  D  �  D  �    �    �  D  �      F  , ,  D  �  D  �    �    �  D  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  D  t  D  <    <    t  D  t      F  , ,  D  t  D  <    <    t  D  t      F  , ,  �  t  �  <  �  <  �  t  �  t      F  , ,  �  t  �  <  �  <  �  t  �  t      F  , ,  $  	�  $  
�  �  
�  �  	�  $  	�      F  , ,  $  	�  $  
�  �  
�  �  	�  $  	�      F  , ,  �  	�  �  
�  |  
�  |  	�  �  	�      F  , ,  �  	�  �  
�  |  
�  |  	�  �  	�      F  , ,  D  	�  D  
�    
�    	�  D  	�      F  , ,  D  	�  D  
�    
�    	�  D  	�      F  , ,  �  �  �  l  |  l  |  �  �  �      F  , ,  �  �  �  l  |  l  |  �  �  �      F  , ,  D  �  D  l    l    �  D  �      F  , ,  D  �  D  l    l    �  D  �      F  , ,  �  �  �  l  �  l  �  �  �  �      F  , ,  �  �  �  l  �  l  �  �  �  �      F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  �  �  �    �        F  , ,  $  �  $  L  �  L  �  �  $  �      F  , ,  $  �  $  L  �  L  �  �  $  �      F  , ,  �  �  �  L  |  L  |  �  �  �      F  , ,  �  �  �  L  |  L  |  �  �  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  $    $  �  �  �  �    $        F  , ,  $    $  �  �  �  �    $        F  , ,  �    �  �  |  �  |    �        F  , ,  �    �  �  |  �  |    �        F  , ,  D    D  �    �      D        F  , ,  D    D  �    �      D        F  , ,  $  �  $  l  �  l  �  �  $  �      F  , ,  $  �  $  l  �  l  �  �  $  �      F  , ,  D  �  D  L    L    �  D  �      F  , ,  D  �  D  L    L    �  D  �      F  , ,  �  �  �  l   l  l   l  �  �  �      F  , ,  �  �  �  l   l  l   l  �  �  �      F  , ,  �  �  �  L   l  L   l  �  �  �      F  , ,  �  �  �  L   l  L   l  �  �  �      F  , ,    �    L  �  L  �  �    �      F  , ,    �    L  �  L  �  �    �      F  , ,  �  �  �  l  �  l  �  �  �  �      F  , ,  �  �  �  l  �  l  �  �  �  �      F  , ,  �  �  �  l  L  l  L  �  �  �      F  , ,  �  �  �  l  L  l  L  �  �  �      F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  L  �  L    �        F  , ,  �    �  �  L  �  L    �        F  , ,  �  �  �  L  L  L  L  �  �  �      F  , ,  �  �  �  L  L  L  L  �  �  �      F  , ,        �  �  �  �            F  , ,        �  �  �  �            F  , ,  �    �  �   l  �   l    �        F  , ,  �    �  �   l  �   l    �        F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,    �    l  �  l  �  �    �      F  , ,    �    l  �  l  �  �    �      F  , ,  "�    "�  �  #�  �  #�    "�        F  , ,  "�    "�  �  #�  �  #�    "�        F  , ,  $T    $T  �  %  �  %    $T        F  , ,  $T    $T  �  %  �  %    $T        F  , ,  %�    %�  �  &�  �  &�    %�        F  , ,  %�    %�  �  &�  �  &�    %�        F  , ,  't    't  �  (<  �  (<    't        F  , ,  't    't  �  (<  �  (<    't        F  , ,  )    )  �  )�  �  )�    )        F  , ,  )    )  �  )�  �  )�    )        F  , ,  *�    *�  �  +\  �  +\    *�        F  , ,  *�    *�  �  +\  �  +\    *�        F  , ,  ,$    ,$  �  ,�  �  ,�    ,$        F  , ,  ,$    ,$  �  ,�  �  ,�    ,$        F  , ,  -�    -�  �  .|  �  .|    -�        F  , ,  -�    -�  �  .|  �  .|    -�        F  , ,  /D    /D  �  0  �  0    /D        F  , ,  /D    /D  �  0  �  0    /D        F  , ,  0�    0�  �  1�  �  1�    0�        F  , ,  0�    0�  �  1�  �  1�    0�        F  , ,  2d    2d  �  3,  �  3,    2d        F  , ,  2d    2d  �  3,  �  3,    2d        F  , ,  3�    3�  �  4�  �  4�    3�        F  , ,  3�    3�  �  4�  �  4�    3�        F  , ,  5�    5�  �  6L  �  6L    5�        F  , ,  5�    5�  �  6L  �  6L    5�        F  , ,  7    7  �  7�  �  7�    7        F  , ,  7    7  �  7�  �  7�    7        F  , ,  8�    8�  �  9l  �  9l    8�        F  , ,  8�    8�  �  9l  �  9l    8�        F  , ,  :4    :4  �  :�  �  :�    :4        F  , ,  :4    :4  �  :�  �  :�    :4        F  , ,  ?    ?  �  ?�  �  ?�    ?        F  , ,  ?    ?  �  ?�  �  ?�    ?        F  , ,  :4  d  :4  ,  :�  ,  :�  d  :4  d      F  , ,  :4  d  :4  ,  :�  ,  :�  d  :4  d      F  , ,  8�  �  8�  �  9l  �  9l  �  8�  �      F  , ,  8�  �  8�  �  9l  �  9l  �  8�  �      F  , ,  :4  �  :4  �  :�  �  :�  �  :4  �      F  , ,  :4  �  :4  �  :�  �  :�  �  :4  �      F  , ,  8�  �  8�  �  9l  �  9l  �  8�  �      F  , ,  8�  �  8�  �  9l  �  9l  �  8�  �      F  , ,  :4  �  :4  �  :�  �  :�  �  :4  �      F  , ,  :4  �  :4  �  :�  �  :�  �  :4  �      F  , ,  8�  �  8�  L  9l  L  9l  �  8�  �      F  , ,  8�  �  8�  L  9l  L  9l  �  8�  �      F  , ,  :4  �  :4  L  :�  L  :�  �  :4  �      F  , ,  :4  �  :4  L  :�  L  :�  �  :4  �      F  , ,  8�    8�  �  9l  �  9l    8�        F  , ,  8�    8�  �  9l  �  9l    8�        F  , ,  :4    :4  �  :�  �  :�    :4        F  , ,  :4    :4  �  :�  �  :�    :4        F  , ,  8�  d  8�  ,  9l  ,  9l  d  8�  d      F  , ,  8�  d  8�  ,  9l  ,  9l  d  8�  d      F  , ,  ?  �  ?  d  ?�  d  ?�  �  ?  �      F  , ,  ?  �  ?  d  ?�  d  ?�  �  ?  �      F  , ,  ?  ,  ?  �  ?�  �  ?�  ,  ?  ,      F  , ,  ?  ,  ?  �  ?�  �  ?�  ,  ?  ,      F  , ,  ?  �  ?  �  ?�  �  ?�  �  ?  �      F  , ,  ?  �  ?  �  ?�  �  ?�  �  ?  �      F  , ,  ?  L  ?    ?�    ?�  L  ?  L      F  , ,  ?  L  ?    ?�    ?�  L  ?  L      F  , ,  7  d  7  ,  7�  ,  7�  d  7  d      F  , ,  7  d  7  ,  7�  ,  7�  d  7  d      F  , ,  3�  d  3�  ,  4�  ,  4�  d  3�  d      F  , ,  3�  d  3�  ,  4�  ,  4�  d  3�  d      F  , ,  5�  d  5�  ,  6L  ,  6L  d  5�  d      F  , ,  5�  d  5�  ,  6L  ,  6L  d  5�  d      F  , ,  0�  �  0�  �  1�  �  1�  �  0�  �      F  , ,  0�  �  0�  �  1�  �  1�  �  0�  �      F  , ,  0�  d  0�  ,  1�  ,  1�  d  0�  d      F  , ,  0�  d  0�  ,  1�  ,  1�  d  0�  d      F  , ,  2d  d  2d  ,  3,  ,  3,  d  2d  d      F  , ,  2d  d  2d  ,  3,  ,  3,  d  2d  d      F  , ,  0�  �  0�  L  1�  L  1�  �  0�  �      F  , ,  0�  �  0�  L  1�  L  1�  �  0�  �      F  , ,  2d  �  2d  L  3,  L  3,  �  2d  �      F  , ,  2d  �  2d  L  3,  L  3,  �  2d  �      F  , ,  3�  �  3�  L  4�  L  4�  �  3�  �      F  , ,  3�  �  3�  L  4�  L  4�  �  3�  �      F  , ,  5�  �  5�  L  6L  L  6L  �  5�  �      F  , ,  5�  �  5�  L  6L  L  6L  �  5�  �      F  , ,  7  �  7  L  7�  L  7�  �  7  �      F  , ,  7  �  7  L  7�  L  7�  �  7  �      F  , ,  2d  �  2d  �  3,  �  3,  �  2d  �      F  , ,  2d  �  2d  �  3,  �  3,  �  2d  �      F  , ,  3�  �  3�  �  4�  �  4�  �  3�  �      F  , ,  3�  �  3�  �  4�  �  4�  �  3�  �      F  , ,  0�    0�  �  1�  �  1�    0�        F  , ,  0�    0�  �  1�  �  1�    0�        F  , ,  2d    2d  �  3,  �  3,    2d        F  , ,  2d    2d  �  3,  �  3,    2d        F  , ,  3�    3�  �  4�  �  4�    3�        F  , ,  3�    3�  �  4�  �  4�    3�        F  , ,  5�    5�  �  6L  �  6L    5�        F  , ,  5�    5�  �  6L  �  6L    5�        F  , ,  7    7  �  7�  �  7�    7        F  , ,  7    7  �  7�  �  7�    7        F  , ,  5�  �  5�  �  6L  �  6L  �  5�  �      F  , ,  5�  �  5�  �  6L  �  6L  �  5�  �      F  , ,  7  �  7  �  7�  �  7�  �  7  �      F  , ,  7  �  7  �  7�  �  7�  �  7  �      F  , ,  0�  �  0�  �  1�  �  1�  �  0�  �      F  , ,  0�  �  0�  �  1�  �  1�  �  0�  �      F  , ,  2d  �  2d  �  3,  �  3,  �  2d  �      F  , ,  2d  �  2d  �  3,  �  3,  �  2d  �      F  , ,  3�  �  3�  �  4�  �  4�  �  3�  �      F  , ,  3�  �  3�  �  4�  �  4�  �  3�  �      F  , ,  5�  �  5�  �  6L  �  6L  �  5�  �      F  , ,  5�  �  5�  �  6L  �  6L  �  5�  �      F  , ,  7  �  7  �  7�  �  7�  �  7  �      F  , ,  7  �  7  �  7�  �  7�  �  7  �      F  , ,  0�  D  0�    1�    1�  D  0�  D      F  , ,  0�  D  0�    1�    1�  D  0�  D      F  , ,  2d  D  2d    3,    3,  D  2d  D      F  , ,  2d  D  2d    3,    3,  D  2d  D      F  , ,  3�  D  3�    4�    4�  D  3�  D      F  , ,  3�  D  3�    4�    4�  D  3�  D      F  , ,  0�  �  0�  \  1�  \  1�  �  0�  �      F  , ,  0�  �  0�  \  1�  \  1�  �  0�  �      F  , ,  2d  �  2d  \  3,  \  3,  �  2d  �      F  , ,  2d  �  2d  \  3,  \  3,  �  2d  �      F  , ,  0�  $  0�  �  1�  �  1�  $  0�  $      F  , ,  0�  $  0�  �  1�  �  1�  $  0�  $      F  , ,  2d  $  2d  �  3,  �  3,  $  2d  $      F  , ,  2d  $  2d  �  3,  �  3,  $  2d  $      F  , ,  3�  $  3�  �  4�  �  4�  $  3�  $      F  , ,  3�  $  3�  �  4�  �  4�  $  3�  $      F  , ,  5�  $  5�  �  6L  �  6L  $  5�  $      F  , ,  5�  $  5�  �  6L  �  6L  $  5�  $      F  , ,  7  $  7  �  7�  �  7�  $  7  $      F  , ,  7  $  7  �  7�  �  7�  $  7  $      F  , ,  0�  �  0�  |  1�  |  1�  �  0�  �      F  , ,  0�  �  0�  |  1�  |  1�  �  0�  �      F  , ,  2d  �  2d  |  3,  |  3,  �  2d  �      F  , ,  2d  �  2d  |  3,  |  3,  �  2d  �      F  , ,  3�  �  3�  |  4�  |  4�  �  3�  �      F  , ,  3�  �  3�  |  4�  |  4�  �  3�  �      F  , ,  5�  �  5�  |  6L  |  6L  �  5�  �      F  , ,  5�  �  5�  |  6L  |  6L  �  5�  �      F  , ,  7  �  7  |  7�  |  7�  �  7  �      F  , ,  7  �  7  |  7�  |  7�  �  7  �      F  , ,  3�  �  3�  \  4�  \  4�  �  3�  �      F  , ,  3�  �  3�  \  4�  \  4�  �  3�  �      F  , ,  5�  �  5�  \  6L  \  6L  �  5�  �      F  , ,  5�  �  5�  \  6L  \  6L  �  5�  �      F  , ,  7  �  7  \  7�  \  7�  �  7  �      F  , ,  7  �  7  \  7�  \  7�  �  7  �      F  , ,  5�  D  5�    6L    6L  D  5�  D      F  , ,  5�  D  5�    6L    6L  D  5�  D      F  , ,  7  D  7    7�    7�  D  7  D      F  , ,  7  D  7    7�    7�  D  7  D      F  , ,  8�  $  8�  �  9l  �  9l  $  8�  $      F  , ,  8�  $  8�  �  9l  �  9l  $  8�  $      F  , ,  8�  �  8�  |  9l  |  9l  �  8�  �      F  , ,  8�  �  8�  |  9l  |  9l  �  8�  �      F  , ,  :4  �  :4  |  :�  |  :�  �  :4  �      F  , ,  :4  �  :4  |  :�  |  :�  �  :4  �      F  , ,  ?  �  ?  �  ?�  �  ?�  �  ?  �      F  , ,  ?  �  ?  �  ?�  �  ?�  �  ?  �      F  , ,  ?  \  ?  $  ?�  $  ?�  \  ?  \      F  , ,  ?  \  ?  $  ?�  $  ?�  \  ?  \      F  , ,  ?  �  ?  �  ?�  �  ?�  �  ?  �      F  , ,  ?  �  ?  �  ?�  �  ?�  �  ?  �      F  , ,  ?  |  ?  D  ?�  D  ?�  |  ?  |      F  , ,  ?  |  ?  D  ?�  D  ?�  |  ?  |      F  , ,  :4  $  :4  �  :�  �  :�  $  :4  $      F  , ,  :4  $  :4  �  :�  �  :�  $  :4  $      F  , ,  8�  D  8�    9l    9l  D  8�  D      F  , ,  8�  D  8�    9l    9l  D  8�  D      F  , ,  :4  D  :4    :�    :�  D  :4  D      F  , ,  :4  D  :4    :�    :�  D  :4  D      F  , ,  8�  �  8�  \  9l  \  9l  �  8�  �      F  , ,  8�  �  8�  \  9l  \  9l  �  8�  �      F  , ,  :4  �  :4  \  :�  \  :�  �  :4  �      F  , ,  :4  �  :4  \  :�  \  :�  �  :4  �      F  , ,  )  �  )  �  )�  �  )�  �  )  �      F  , ,  )  �  )  �  )�  �  )�  �  )  �      F  , ,  )  �  )  \  )�  \  )�  �  )  �      F  , ,  )  �  )  \  )�  \  )�  �  )  �      F  , ,  )    )  �  )�  �  )�    )        F  , ,  )    )  �  )�  �  )�    )        F  , ,  )  D  )    )�    )�  D  )  D      F  , ,  )  D  )    )�    )�  D  )  D      F  , ,  )  �  )  �  )�  �  )�  �  )  �      F  , ,  )  �  )  �  )�  �  )�  �  )  �      F  , ,  )  $  )  �  )�  �  )�  $  )  $      F  , ,  )  $  )  �  )�  �  )�  $  )  $      F  , ,  )  �  )  |  )�  |  )�  �  )  �      F  , ,  )  �  )  |  )�  |  )�  �  )  �      F  , ,  )  d  )  ,  )�  ,  )�  d  )  d      F  , ,  )  d  )  ,  )�  ,  )�  d  )  d      F  , ,  )  �  )  L  )�  L  )�  �  )  �      F  , ,  )  �  )  L  )�  L  )�  �  )  �      F  , ,  ,$    ,$  �  ,�  �  ,�    ,$        F  , ,  ,$    ,$  �  ,�  �  ,�    ,$        F  , ,  -�    -�  �  .|  �  .|    -�        F  , ,  -�    -�  �  .|  �  .|    -�        F  , ,  /D    /D  �  0  �  0    /D        F  , ,  /D    /D  �  0  �  0    /D        F  , ,  ,$  �  ,$  �  ,�  �  ,�  �  ,$  �      F  , ,  ,$  �  ,$  �  ,�  �  ,�  �  ,$  �      F  , ,  -�  �  -�  �  .|  �  .|  �  -�  �      F  , ,  -�  �  -�  �  .|  �  .|  �  -�  �      F  , ,  /D  �  /D  L  0  L  0  �  /D  �      F  , ,  /D  �  /D  L  0  L  0  �  /D  �      F  , ,  *�  �  *�  �  +\  �  +\  �  *�  �      F  , ,  *�  �  *�  �  +\  �  +\  �  *�  �      F  , ,  ,$  �  ,$  �  ,�  �  ,�  �  ,$  �      F  , ,  ,$  �  ,$  �  ,�  �  ,�  �  ,$  �      F  , ,  -�  �  -�  �  .|  �  .|  �  -�  �      F  , ,  -�  �  -�  �  .|  �  .|  �  -�  �      F  , ,  /D  �  /D  �  0  �  0  �  /D  �      F  , ,  /D  �  /D  �  0  �  0  �  /D  �      F  , ,  /D  �  /D  �  0  �  0  �  /D  �      F  , ,  /D  �  /D  �  0  �  0  �  /D  �      F  , ,  *�  �  *�  �  +\  �  +\  �  *�  �      F  , ,  *�  �  *�  �  +\  �  +\  �  *�  �      F  , ,  *�  d  *�  ,  +\  ,  +\  d  *�  d      F  , ,  *�  d  *�  ,  +\  ,  +\  d  *�  d      F  , ,  ,$  d  ,$  ,  ,�  ,  ,�  d  ,$  d      F  , ,  ,$  d  ,$  ,  ,�  ,  ,�  d  ,$  d      F  , ,  -�  d  -�  ,  .|  ,  .|  d  -�  d      F  , ,  -�  d  -�  ,  .|  ,  .|  d  -�  d      F  , ,  /D  d  /D  ,  0  ,  0  d  /D  d      F  , ,  /D  d  /D  ,  0  ,  0  d  /D  d      F  , ,  *�    *�  �  +\  �  +\    *�        F  , ,  *�    *�  �  +\  �  +\    *�        F  , ,  *�  �  *�  L  +\  L  +\  �  *�  �      F  , ,  *�  �  *�  L  +\  L  +\  �  *�  �      F  , ,  ,$  �  ,$  L  ,�  L  ,�  �  ,$  �      F  , ,  ,$  �  ,$  L  ,�  L  ,�  �  ,$  �      F  , ,  -�  �  -�  L  .|  L  .|  �  -�  �      F  , ,  -�  �  -�  L  .|  L  .|  �  -�  �      F  , ,  "�    "�  �  #�  �  #�    "�        F  , ,  "�    "�  �  #�  �  #�    "�        F  , ,  $T    $T  �  %  �  %    $T        F  , ,  $T    $T  �  %  �  %    $T        F  , ,  $T  d  $T  ,  %  ,  %  d  $T  d      F  , ,  $T  d  $T  ,  %  ,  %  d  $T  d      F  , ,  %�  d  %�  ,  &�  ,  &�  d  %�  d      F  , ,  %�  d  %�  ,  &�  ,  &�  d  %�  d      F  , ,  't  d  't  ,  (<  ,  (<  d  't  d      F  , ,  't  d  't  ,  (<  ,  (<  d  't  d      F  , ,  %�    %�  �  &�  �  &�    %�        F  , ,  %�    %�  �  &�  �  &�    %�        F  , ,  "�  d  "�  ,  #�  ,  #�  d  "�  d      F  , ,  "�  d  "�  ,  #�  ,  #�  d  "�  d      F  , ,  "�  �  "�  �  #�  �  #�  �  "�  �      F  , ,  "�  �  "�  �  #�  �  #�  �  "�  �      F  , ,  $T  �  $T  �  %  �  %  �  $T  �      F  , ,  $T  �  $T  �  %  �  %  �  $T  �      F  , ,  %�  �  %�  �  &�  �  &�  �  %�  �      F  , ,  %�  �  %�  �  &�  �  &�  �  %�  �      F  , ,  't  �  't  �  (<  �  (<  �  't  �      F  , ,  't  �  't  �  (<  �  (<  �  't  �      F  , ,  "�  �  "�  �  #�  �  #�  �  "�  �      F  , ,  "�  �  "�  �  #�  �  #�  �  "�  �      F  , ,  "�  �  "�  L  #�  L  #�  �  "�  �      F  , ,  "�  �  "�  L  #�  L  #�  �  "�  �      F  , ,  $T  �  $T  L  %  L  %  �  $T  �      F  , ,  $T  �  $T  L  %  L  %  �  $T  �      F  , ,  %�  �  %�  L  &�  L  &�  �  %�  �      F  , ,  %�  �  %�  L  &�  L  &�  �  %�  �      F  , ,  't  �  't  L  (<  L  (<  �  't  �      F  , ,  't  �  't  L  (<  L  (<  �  't  �      F  , ,  't    't  �  (<  �  (<    't        F  , ,  't    't  �  (<  �  (<    't        F  , ,  $T  �  $T  �  %  �  %  �  $T  �      F  , ,  $T  �  $T  �  %  �  %  �  $T  �      F  , ,  %�  �  %�  �  &�  �  &�  �  %�  �      F  , ,  %�  �  %�  �  &�  �  &�  �  %�  �      F  , ,  't  �  't  �  (<  �  (<  �  't  �      F  , ,  't  �  't  �  (<  �  (<  �  't  �      F  , ,  't  �  't  |  (<  |  (<  �  't  �      F  , ,  't  �  't  |  (<  |  (<  �  't  �      F  , ,  "�  $  "�  �  #�  �  #�  $  "�  $      F  , ,  "�  $  "�  �  #�  �  #�  $  "�  $      F  , ,  $T  $  $T  �  %  �  %  $  $T  $      F  , ,  $T  $  $T  �  %  �  %  $  $T  $      F  , ,  %�  $  %�  �  &�  �  &�  $  %�  $      F  , ,  %�  $  %�  �  &�  �  &�  $  %�  $      F  , ,  't  $  't  �  (<  �  (<  $  't  $      F  , ,  't  $  't  �  (<  �  (<  $  't  $      F  , ,  %�  �  %�  \  &�  \  &�  �  %�  �      F  , ,  %�  �  %�  \  &�  \  &�  �  %�  �      F  , ,  't  �  't  \  (<  \  (<  �  't  �      F  , ,  't  �  't  \  (<  \  (<  �  't  �      F  , ,  "�  �  "�  \  #�  \  #�  �  "�  �      F  , ,  "�  �  "�  \  #�  \  #�  �  "�  �      F  , ,  $T  �  $T  \  %  \  %  �  $T  �      F  , ,  $T  �  $T  \  %  \  %  �  $T  �      F  , ,  "�  D  "�    #�    #�  D  "�  D      F  , ,  "�  D  "�    #�    #�  D  "�  D      F  , ,  $T  D  $T    %    %  D  $T  D      F  , ,  $T  D  $T    %    %  D  $T  D      F  , ,  %�  D  %�    &�    &�  D  %�  D      F  , ,  %�  D  %�    &�    &�  D  %�  D      F  , ,  't  D  't    (<    (<  D  't  D      F  , ,  't  D  't    (<    (<  D  't  D      F  , ,  "�  �  "�  |  #�  |  #�  �  "�  �      F  , ,  "�  �  "�  |  #�  |  #�  �  "�  �      F  , ,  $T  �  $T  |  %  |  %  �  $T  �      F  , ,  $T  �  $T  |  %  |  %  �  $T  �      F  , ,  %�  �  %�  |  &�  |  &�  �  %�  �      F  , ,  %�  �  %�  |  &�  |  &�  �  %�  �      F  , ,  *�  �  *�  \  +\  \  +\  �  *�  �      F  , ,  *�  �  *�  \  +\  \  +\  �  *�  �      F  , ,  -�  D  -�    .|    .|  D  -�  D      F  , ,  -�  D  -�    .|    .|  D  -�  D      F  , ,  /D  D  /D    0    0  D  /D  D      F  , ,  /D  D  /D    0    0  D  /D  D      F  , ,  ,$  �  ,$  \  ,�  \  ,�  �  ,$  �      F  , ,  ,$  �  ,$  \  ,�  \  ,�  �  ,$  �      F  , ,  *�  $  *�  �  +\  �  +\  $  *�  $      F  , ,  *�  $  *�  �  +\  �  +\  $  *�  $      F  , ,  *�  D  *�    +\    +\  D  *�  D      F  , ,  *�  D  *�    +\    +\  D  *�  D      F  , ,  ,$  D  ,$    ,�    ,�  D  ,$  D      F  , ,  ,$  D  ,$    ,�    ,�  D  ,$  D      F  , ,  ,$  $  ,$  �  ,�  �  ,�  $  ,$  $      F  , ,  ,$  $  ,$  �  ,�  �  ,�  $  ,$  $      F  , ,  -�  $  -�  �  .|  �  .|  $  -�  $      F  , ,  -�  $  -�  �  .|  �  .|  $  -�  $      F  , ,  /D  $  /D  �  0  �  0  $  /D  $      F  , ,  /D  $  /D  �  0  �  0  $  /D  $      F  , ,  -�  �  -�  \  .|  \  .|  �  -�  �      F  , ,  -�  �  -�  \  .|  \  .|  �  -�  �      F  , ,  /D  �  /D  \  0  \  0  �  /D  �      F  , ,  /D  �  /D  \  0  \  0  �  /D  �      F  , ,  *�  �  *�  |  +\  |  +\  �  *�  �      F  , ,  *�  �  *�  |  +\  |  +\  �  *�  �      F  , ,  ,$  �  ,$  |  ,�  |  ,�  �  ,$  �      F  , ,  ,$  �  ,$  |  ,�  |  ,�  �  ,$  �      F  , ,  -�  �  -�  |  .|  |  .|  �  -�  �      F  , ,  -�  �  -�  |  .|  |  .|  �  -�  �      F  , ,  /D  �  /D  |  0  |  0  �  /D  �      F  , ,  /D  �  /D  |  0  |  0  �  /D  �      F  , ,  )  T  )    )�    )�  T  )  T      F  , ,  )  T  )    )�    )�  T  )  T      F  , ,  )  �  )  L  )�  L  )�  �  )  �      F  , ,  )  �  )  L  )�  L  )�  �  )  �      F  , ,  )  	�  )  
�  )�  
�  )�  	�  )  	�      F  , ,  )  	�  )  
�  )�  
�  )�  	�  )  	�      F  , ,  )  t  )  <  )�  <  )�  t  )  t      F  , ,  )  t  )  <  )�  <  )�  t  )  t      F  , ,  "�  4  "�  �  #�  �  #�  4  "�  4      F  , ,  "�  4  "�  �  #�  �  #�  4  "�  4      F  , ,  $T  4  $T  �  %  �  %  4  $T  4      F  , ,  $T  4  $T  �  %  �  %  4  $T  4      F  , ,  %�  4  %�  �  &�  �  &�  4  %�  4      F  , ,  %�  4  %�  �  &�  �  &�  4  %�  4      F  , ,  't  4  't  �  (<  �  (<  4  't  4      F  , ,  't  4  't  �  (<  �  (<  4  't  4      F  , ,  )  4  )  �  )�  �  )�  4  )  4      F  , ,  )  4  )  �  )�  �  )�  4  )  4      F  , ,  *�  4  *�  �  +\  �  +\  4  *�  4      F  , ,  *�  4  *�  �  +\  �  +\  4  *�  4      F  , ,  ,$  4  ,$  �  ,�  �  ,�  4  ,$  4      F  , ,  ,$  4  ,$  �  ,�  �  ,�  4  ,$  4      F  , ,  -�  4  -�  �  .|  �  .|  4  -�  4      F  , ,  -�  4  -�  �  .|  �  .|  4  -�  4      F  , ,  /D  4  /D  �  0  �  0  4  /D  4      F  , ,  /D  4  /D  �  0  �  0  4  /D  4      F  , ,  )    )  �  )�  �  )�    )        F  , ,  )    )  �  )�  �  )�    )        F  , ,  )  �  )  l  )�  l  )�  �  )  �      F  , ,  )  �  )  l  )�  l  )�  �  )  �      F  , ,  )  �  )  �  )�  �  )�  �  )  �      F  , ,  )  �  )  �  )�  �  )�  �  )  �      F  , ,  ,$  T  ,$    ,�    ,�  T  ,$  T      F  , ,  ,$  T  ,$    ,�    ,�  T  ,$  T      F  , ,  *�  	�  *�  
�  +\  
�  +\  	�  *�  	�      F  , ,  *�  	�  *�  
�  +\  
�  +\  	�  *�  	�      F  , ,  ,$  	�  ,$  
�  ,�  
�  ,�  	�  ,$  	�      F  , ,  ,$  	�  ,$  
�  ,�  
�  ,�  	�  ,$  	�      F  , ,  -�  	�  -�  
�  .|  
�  .|  	�  -�  	�      F  , ,  -�  	�  -�  
�  .|  
�  .|  	�  -�  	�      F  , ,  -�  T  -�    .|    .|  T  -�  T      F  , ,  -�  T  -�    .|    .|  T  -�  T      F  , ,  *�  t  *�  <  +\  <  +\  t  *�  t      F  , ,  *�  t  *�  <  +\  <  +\  t  *�  t      F  , ,  ,$  t  ,$  <  ,�  <  ,�  t  ,$  t      F  , ,  ,$  t  ,$  <  ,�  <  ,�  t  ,$  t      F  , ,  -�  t  -�  <  .|  <  .|  t  -�  t      F  , ,  -�  t  -�  <  .|  <  .|  t  -�  t      F  , ,  /D  	�  /D  
�  0  
�  0  	�  /D  	�      F  , ,  /D  	�  /D  
�  0  
�  0  	�  /D  	�      F  , ,  /D  t  /D  <  0  <  0  t  /D  t      F  , ,  /D  t  /D  <  0  <  0  t  /D  t      F  , ,  /D  T  /D    0    0  T  /D  T      F  , ,  /D  T  /D    0    0  T  /D  T      F  , ,  *�  T  *�    +\    +\  T  *�  T      F  , ,  *�  T  *�    +\    +\  T  *�  T      F  , ,  *�  �  *�  �  +\  �  +\  �  *�  �      F  , ,  *�  �  *�  �  +\  �  +\  �  *�  �      F  , ,  ,$  �  ,$  �  ,�  �  ,�  �  ,$  �      F  , ,  ,$  �  ,$  �  ,�  �  ,�  �  ,$  �      F  , ,  -�  �  -�  �  .|  �  .|  �  -�  �      F  , ,  -�  �  -�  �  .|  �  .|  �  -�  �      F  , ,  /D  �  /D  �  0  �  0  �  /D  �      F  , ,  /D  �  /D  �  0  �  0  �  /D  �      F  , ,  %�  �  %�  �  &�  �  &�  �  %�  �      F  , ,  %�  �  %�  �  &�  �  &�  �  %�  �      F  , ,  't  �  't  �  (<  �  (<  �  't  �      F  , ,  't  �  't  �  (<  �  (<  �  't  �      F  , ,  "�  	�  "�  
�  #�  
�  #�  	�  "�  	�      F  , ,  "�  	�  "�  
�  #�  
�  #�  	�  "�  	�      F  , ,  $T  	�  $T  
�  %  
�  %  	�  $T  	�      F  , ,  $T  	�  $T  
�  %  
�  %  	�  $T  	�      F  , ,  "�  t  "�  <  #�  <  #�  t  "�  t      F  , ,  "�  t  "�  <  #�  <  #�  t  "�  t      F  , ,  $T  t  $T  <  %  <  %  t  $T  t      F  , ,  $T  t  $T  <  %  <  %  t  $T  t      F  , ,  %�  t  %�  <  &�  <  &�  t  %�  t      F  , ,  %�  t  %�  <  &�  <  &�  t  %�  t      F  , ,  't  t  't  <  (<  <  (<  t  't  t      F  , ,  't  t  't  <  (<  <  (<  t  't  t      F  , ,  %�  	�  %�  
�  &�  
�  &�  	�  %�  	�      F  , ,  %�  	�  %�  
�  &�  
�  &�  	�  %�  	�      F  , ,  't  	�  't  
�  (<  
�  (<  	�  't  	�      F  , ,  't  	�  't  
�  (<  
�  (<  	�  't  	�      F  , ,  "�  T  "�    #�    #�  T  "�  T      F  , ,  "�  T  "�    #�    #�  T  "�  T      F  , ,  $T  T  $T    %    %  T  $T  T      F  , ,  $T  T  $T    %    %  T  $T  T      F  , ,  %�  T  %�    &�    &�  T  %�  T      F  , ,  %�  T  %�    &�    &�  T  %�  T      F  , ,  't  T  't    (<    (<  T  't  T      F  , ,  't  T  't    (<    (<  T  't  T      F  , ,  "�  �  "�  �  #�  �  #�  �  "�  �      F  , ,  "�  �  "�  �  #�  �  #�  �  "�  �      F  , ,  $T  �  $T  �  %  �  %  �  $T  �      F  , ,  $T  �  $T  �  %  �  %  �  $T  �      F  , ,  %�  �  %�  L  &�  L  &�  �  %�  �      F  , ,  %�  �  %�  L  &�  L  &�  �  %�  �      F  , ,  't  �  't  L  (<  L  (<  �  't  �      F  , ,  't  �  't  L  (<  L  (<  �  't  �      F  , ,  "�    "�  �  #�  �  #�    "�        F  , ,  "�    "�  �  #�  �  #�    "�        F  , ,  $T    $T  �  %  �  %    $T        F  , ,  $T    $T  �  %  �  %    $T        F  , ,  %�    %�  �  &�  �  &�    %�        F  , ,  %�    %�  �  &�  �  &�    %�        F  , ,  't    't  �  (<  �  (<    't        F  , ,  't    't  �  (<  �  (<    't        F  , ,  "�  �  "�  l  #�  l  #�  �  "�  �      F  , ,  "�  �  "�  l  #�  l  #�  �  "�  �      F  , ,  $T  �  $T  l  %  l  %  �  $T  �      F  , ,  $T  �  $T  l  %  l  %  �  $T  �      F  , ,  %�  �  %�  l  &�  l  &�  �  %�  �      F  , ,  %�  �  %�  l  &�  l  &�  �  %�  �      F  , ,  "�  �  "�  L  #�  L  #�  �  "�  �      F  , ,  "�  �  "�  L  #�  L  #�  �  "�  �      F  , ,  't  �  't  l  (<  l  (<  �  't  �      F  , ,  't  �  't  l  (<  l  (<  �  't  �      F  , ,  $T  �  $T  L  %  L  %  �  $T  �      F  , ,  $T  �  $T  L  %  L  %  �  $T  �      F  , ,  *�  �  *�  L  +\  L  +\  �  *�  �      F  , ,  *�  �  *�  L  +\  L  +\  �  *�  �      F  , ,  /D  �  /D  L  0  L  0  �  /D  �      F  , ,  /D  �  /D  L  0  L  0  �  /D  �      F  , ,  ,$  �  ,$  L  ,�  L  ,�  �  ,$  �      F  , ,  ,$  �  ,$  L  ,�  L  ,�  �  ,$  �      F  , ,  -�  �  -�  L  .|  L  .|  �  -�  �      F  , ,  -�  �  -�  L  .|  L  .|  �  -�  �      F  , ,  /D  �  /D  l  0  l  0  �  /D  �      F  , ,  /D  �  /D  l  0  l  0  �  /D  �      F  , ,  *�  �  *�  l  +\  l  +\  �  *�  �      F  , ,  *�  �  *�  l  +\  l  +\  �  *�  �      F  , ,  *�    *�  �  +\  �  +\    *�        F  , ,  *�    *�  �  +\  �  +\    *�        F  , ,  ,$    ,$  �  ,�  �  ,�    ,$        F  , ,  ,$    ,$  �  ,�  �  ,�    ,$        F  , ,  -�    -�  �  .|  �  .|    -�        F  , ,  -�    -�  �  .|  �  .|    -�        F  , ,  /D    /D  �  0  �  0    /D        F  , ,  /D    /D  �  0  �  0    /D        F  , ,  ,$  �  ,$  l  ,�  l  ,�  �  ,$  �      F  , ,  ,$  �  ,$  l  ,�  l  ,�  �  ,$  �      F  , ,  -�  �  -�  l  .|  l  .|  �  -�  �      F  , ,  -�  �  -�  l  .|  l  .|  �  -�  �      F  , ,  0�  4  0�  �  1�  �  1�  4  0�  4      F  , ,  0�  4  0�  �  1�  �  1�  4  0�  4      F  , ,  2d  4  2d  �  3,  �  3,  4  2d  4      F  , ,  2d  4  2d  �  3,  �  3,  4  2d  4      F  , ,  3�  4  3�  �  4�  �  4�  4  3�  4      F  , ,  3�  4  3�  �  4�  �  4�  4  3�  4      F  , ,  5�  4  5�  �  6L  �  6L  4  5�  4      F  , ,  5�  4  5�  �  6L  �  6L  4  5�  4      F  , ,  7  4  7  �  7�  �  7�  4  7  4      F  , ,  7  4  7  �  7�  �  7�  4  7  4      F  , ,  8�  4  8�  �  9l  �  9l  4  8�  4      F  , ,  8�  4  8�  �  9l  �  9l  4  8�  4      F  , ,  :4  4  :4  �  :�  �  :�  4  :4  4      F  , ,  :4  4  :4  �  :�  �  :�  4  :4  4      F  , ,  ?  �  ?  	�  ?�  	�  ?�  �  ?  �      F  , ,  ?  �  ?  	�  ?�  	�  ?�  �  ?  �      F  , ,  ?  
�  ?  T  ?�  T  ?�  
�  ?  
�      F  , ,  ?  
�  ?  T  ?�  T  ?�  
�  ?  
�      F  , ,  ?    ?  �  ?�  �  ?�    ?        F  , ,  ?    ?  �  ?�  �  ?�    ?        F  , ,  ?  �  ?  t  ?�  t  ?�  �  ?  �      F  , ,  ?  �  ?  t  ?�  t  ?�  �  ?  �      F  , ,  ?  <  ?    ?�    ?�  <  ?  <      F  , ,  ?  <  ?    ?�    ?�  <  ?  <      F  , ,  :4  t  :4  <  :�  <  :�  t  :4  t      F  , ,  :4  t  :4  <  :�  <  :�  t  :4  t      F  , ,  8�  	�  8�  
�  9l  
�  9l  	�  8�  	�      F  , ,  8�  	�  8�  
�  9l  
�  9l  	�  8�  	�      F  , ,  8�  �  8�  �  9l  �  9l  �  8�  �      F  , ,  8�  �  8�  �  9l  �  9l  �  8�  �      F  , ,  :4  �  :4  �  :�  �  :�  �  :4  �      F  , ,  :4  �  :4  �  :�  �  :�  �  :4  �      F  , ,  :4  	�  :4  
�  :�  
�  :�  	�  :4  	�      F  , ,  :4  	�  :4  
�  :�  
�  :�  	�  :4  	�      F  , ,  8�  T  8�    9l    9l  T  8�  T      F  , ,  8�  T  8�    9l    9l  T  8�  T      F  , ,  :4  T  :4    :�    :�  T  :4  T      F  , ,  :4  T  :4    :�    :�  T  :4  T      F  , ,  8�  t  8�  <  9l  <  9l  t  8�  t      F  , ,  8�  t  8�  <  9l  <  9l  t  8�  t      F  , ,  0�  T  0�    1�    1�  T  0�  T      F  , ,  0�  T  0�    1�    1�  T  0�  T      F  , ,  3�  t  3�  <  4�  <  4�  t  3�  t      F  , ,  3�  t  3�  <  4�  <  4�  t  3�  t      F  , ,  0�  t  0�  <  1�  <  1�  t  0�  t      F  , ,  0�  t  0�  <  1�  <  1�  t  0�  t      F  , ,  0�  	�  0�  
�  1�  
�  1�  	�  0�  	�      F  , ,  0�  	�  0�  
�  1�  
�  1�  	�  0�  	�      F  , ,  2d  	�  2d  
�  3,  
�  3,  	�  2d  	�      F  , ,  2d  	�  2d  
�  3,  
�  3,  	�  2d  	�      F  , ,  3�  	�  3�  
�  4�  
�  4�  	�  3�  	�      F  , ,  3�  	�  3�  
�  4�  
�  4�  	�  3�  	�      F  , ,  5�  	�  5�  
�  6L  
�  6L  	�  5�  	�      F  , ,  5�  	�  5�  
�  6L  
�  6L  	�  5�  	�      F  , ,  7  	�  7  
�  7�  
�  7�  	�  7  	�      F  , ,  7  	�  7  
�  7�  
�  7�  	�  7  	�      F  , ,  5�  t  5�  <  6L  <  6L  t  5�  t      F  , ,  5�  t  5�  <  6L  <  6L  t  5�  t      F  , ,  0�  �  0�  �  1�  �  1�  �  0�  �      F  , ,  0�  �  0�  �  1�  �  1�  �  0�  �      F  , ,  2d  �  2d  �  3,  �  3,  �  2d  �      F  , ,  2d  �  2d  �  3,  �  3,  �  2d  �      F  , ,  3�  �  3�  �  4�  �  4�  �  3�  �      F  , ,  3�  �  3�  �  4�  �  4�  �  3�  �      F  , ,  5�  �  5�  �  6L  �  6L  �  5�  �      F  , ,  5�  �  5�  �  6L  �  6L  �  5�  �      F  , ,  7  �  7  �  7�  �  7�  �  7  �      F  , ,  7  �  7  �  7�  �  7�  �  7  �      F  , ,  7  t  7  <  7�  <  7�  t  7  t      F  , ,  7  t  7  <  7�  <  7�  t  7  t      F  , ,  2d  T  2d    3,    3,  T  2d  T      F  , ,  2d  T  2d    3,    3,  T  2d  T      F  , ,  3�  T  3�    4�    4�  T  3�  T      F  , ,  3�  T  3�    4�    4�  T  3�  T      F  , ,  5�  T  5�    6L    6L  T  5�  T      F  , ,  5�  T  5�    6L    6L  T  5�  T      F  , ,  7  T  7    7�    7�  T  7  T      F  , ,  7  T  7    7�    7�  T  7  T      F  , ,  2d  t  2d  <  3,  <  3,  t  2d  t      F  , ,  2d  t  2d  <  3,  <  3,  t  2d  t      F  , ,  7  �  7  l  7�  l  7�  �  7  �      F  , ,  7  �  7  l  7�  l  7�  �  7  �      F  , ,  5�    5�  �  6L  �  6L    5�        F  , ,  5�    5�  �  6L  �  6L    5�        F  , ,  7    7  �  7�  �  7�    7        F  , ,  7    7  �  7�  �  7�    7        F  , ,  0�  �  0�  l  1�  l  1�  �  0�  �      F  , ,  0�  �  0�  l  1�  l  1�  �  0�  �      F  , ,  2d  �  2d  l  3,  l  3,  �  2d  �      F  , ,  2d  �  2d  l  3,  l  3,  �  2d  �      F  , ,  3�  �  3�  l  4�  l  4�  �  3�  �      F  , ,  3�  �  3�  l  4�  l  4�  �  3�  �      F  , ,  0�    0�  �  1�  �  1�    0�        F  , ,  0�    0�  �  1�  �  1�    0�        F  , ,  0�  �  0�  L  1�  L  1�  �  0�  �      F  , ,  0�  �  0�  L  1�  L  1�  �  0�  �      F  , ,  2d  �  2d  L  3,  L  3,  �  2d  �      F  , ,  2d  �  2d  L  3,  L  3,  �  2d  �      F  , ,  3�  �  3�  L  4�  L  4�  �  3�  �      F  , ,  3�  �  3�  L  4�  L  4�  �  3�  �      F  , ,  2d    2d  �  3,  �  3,    2d        F  , ,  2d    2d  �  3,  �  3,    2d        F  , ,  3�    3�  �  4�  �  4�    3�        F  , ,  3�    3�  �  4�  �  4�    3�        F  , ,  5�  �  5�  l  6L  l  6L  �  5�  �      F  , ,  5�  �  5�  l  6L  l  6L  �  5�  �      F  , ,  5�  �  5�  L  6L  L  6L  �  5�  �      F  , ,  5�  �  5�  L  6L  L  6L  �  5�  �      F  , ,  7  �  7  L  7�  L  7�  �  7  �      F  , ,  7  �  7  L  7�  L  7�  �  7  �      F  , ,  ?  �  ?  �  ?�  �  ?�  �  ?  �      F  , ,  ?  �  ?  �  ?�  �  ?�  �  ?  �      F  , ,  ?  L  ?    ?�    ?�  L  ?  L      F  , ,  ?  L  ?    ?�    ?�  L  ?  L      F  , ,  ?  �  ?  �  ?�  �  ?�  �  ?  �      F  , ,  ?  �  ?  �  ?�  �  ?�  �  ?  �      F  , ,  ?  l  ?  4  ?�  4  ?�  l  ?  l      F  , ,  ?  l  ?  4  ?�  4  ?�  l  ?  l      F  , ,  8�  �  8�  l  9l  l  9l  �  8�  �      F  , ,  8�  �  8�  l  9l  l  9l  �  8�  �      F  , ,  :4  �  :4  l  :�  l  :�  �  :4  �      F  , ,  :4  �  :4  l  :�  l  :�  �  :4  �      F  , ,  8�    8�  �  9l  �  9l    8�        F  , ,  8�    8�  �  9l  �  9l    8�        F  , ,  :4    :4  �  :�  �  :�    :4        F  , ,  :4    :4  �  :�  �  :�    :4        F  , ,  ?  ,  ?  �  ?�  �  ?�  ,  ?  ,      F  , ,  ?  ,  ?  �  ?�  �  ?�  ,  ?  ,      F  , ,  8�  �  8�  L  9l  L  9l  �  8�  �      F  , ,  8�  �  8�  L  9l  L  9l  �  8�  �      F  , ,  :4  �  :4  L  :�  L  :�  �  :4  �      F  , ,  :4  �  :4  L  :�  L  :�  �  :4  �      �   ,              >�  >�  >�  >�                  Y  , ,  �  �  �  <�  <�  <�  <�  �  �  �     �     0�     0 *sky130_fd_pr__res_high_po_0p35_8WX6FW    �     0�     0 *sky130_fd_pr__res_high_po_0p35_ZNVMZH    �     0�     0 *sky130_fd_pr__res_high_po_0p35_TFWMD7    �     0�     0 *sky130_fd_pr__res_high_po_0p35_EN8PRN    �     0�     0 *sky130_fd_pr__res_xhigh_po_0p35_CJJ24B   �     0�     0 via_new$1  	   D   !     �           �       	   E   !     �           �       	   F   !     �           �       	   G   !     �           �          D  , ,   �����   �   K  '   K  '����   �����      D  , ,  �����  �   K  g   K  g����  �����      D  , ,  ����     K  �   K  �����  ����      D  , ,  Q����  Q   K  �   K  �����  Q����      D  , ,  �����  �   K  '   K  '����  �����      D  , ,  �����  �   K  g   K  g����  �����      D  , ,  ����     K  �   K  �����  ����      D  , ,  	Q����  	Q   K  	�   K  	�����  	Q����      D  , ,  
�����  
�   K  '   K  '����  
�����      E  , ,   �����   �   d  �   d  �����   �����      E  , ,  X����  X   d      d   ����  X����      E  , ,  �����  �   d  �   d  �����  �����      E  , ,  x����  x   d  @   d  @����  x����      E  , ,  ����     d  �   d  �����  ����      E  , ,  �����  �   d  	`   d  	`����  �����      E  , ,  
(����  
(   d  
�   d  
�����  
(����      F  , ,   �����   �   d  �   d  �����   �����      F  , ,  X����  X   d      d   ����  X����      F  , ,  �����  �   d  �   d  �����  �����      F  , ,  x����  x   d  @   d  @����  x����      F  , ,  ����     d  �   d  �����  ����      F  , ,  �����  �   d  	`   d  	`����  �����      F  , ,  
(����  
(   d  
�   d  
�����  
(����     �     0�     0 *sky130_fd_pr__res_high_po_0p35_LCRD8L     B   ,��f��{X��f��|���0���|���0���{X��f��{X      B   ,��f������f������0�������0�������f����      B   ,��f������f���"��0����"��0�������f����      _   ,����z�����}��0���}��0���z�����z�      _   ,�����/�����K��0����K��0����/�����/      _   ,�����e��������0�������0����e�����e      C   ,�����x��������������������x������x�      C   ,�����x������yx��2~��yx��2~��x������x�      C   ,��f��{X��f��|������|������{X��f��{X      C   ,��f������f��������������������f����      C   ,��f������f���"������"���������f����      C   ,��(.��{X��(.��|���0���|���0���{X��(.��{X      C   ,��(.������(.������0�������0�������(.����      C   ,��(.������(.���"��0����"��0�������(.����      C   ,���������������2~������2~���������      C   ,��2~��x���2~������3(������3(��x���2~��x�      D   ,�����{������|������|������{������{�      D   ,�����������������������������������      D   ,�����������������������������������      D   ,��(G��{���(G��|���0���|���0���{���(G��{�      D   ,��(G������(G������0�������0�������(G����      D   ,��(G������(G������0�������0�������(G����      C  , ,�����{������|\��t��|\��t��{������{�      C  , ,����������������t������t�����������      C  , ,���������������t������t���������      C  , ,��2��{���2��|\�����|\�����{���2��{�      C  , ,��2������2��������������������2����      C  , ,��2�����2�������������������2���      C  , ,�����{������|\��D��|\��D��{������{�      C  , ,����������������D������D�����������      C  , ,���������������D������D���������      C  , ,��	��{���	��|\��	���|\��	���{���	��{�      C  , ,��	������	������	�������	�������	����      C  , ,��	�����	������	�������	������	���      C  , ,��
j��{���
j��|\����|\����{���
j��{�      C  , ,��
j������
j������������������
j����      C  , ,��
j�����
j�����������������
j���      C  , ,�����{������|\��|��|\��|��{������{�      C  , ,����������������|������|�����������      C  , ,���������������|������|���������      C  , ,��(���{���(���|\��)7��|\��)7��{���(���{�      C  , ,��(�������(�������)7������)7������(�����      C  , ,��(������(�������)7������)7�����(����      C  , ,��)���{���)���|\��*���|\��*���{���)���{�      C  , ,��)�������)�������*�������*�������)�����      C  , ,��)������)�������*�������*������)����      C  , ,��+]��{���+]��|\��,��|\��,��{���+]��{�      C  , ,��+]������+]������,������,������+]����      C  , ,��+]�����+]������,������,�����+]���      C  , ,��,���{���,���|\��-o��|\��-o��{���,���{�      C  , ,��,�������,�������-o������-o������,�����      C  , ,��,������,�������-o������-o�����,����      C  , ,��.-��{���.-��|\��.���|\��.���{���.-��{�      C  , ,��.-������.-������.�������.�������.-����      C  , ,��.-�����.-������.�������.������.-���      C  , ,��/���{���/���|\��0?��|\��0?��{���/���{�      C  , ,��/�������/�������0?������0?������/�����      C  , ,��/������/�������0?������0?�����/����      ^   ,��_��xQ��_���)�����)����xQ��_��xQ      ^   ,����xQ����}$��2��}$��2��xQ����xQ      ^   ,����� �����Z��2���Z��2��� �����       ^   ,�����V�����)��2���)��2���V�����V      ^   ,��2��xQ��2���)��3����)��3���xQ��2��xQ      A  , ,�����x��������������������x������x�      A  , ,�����x������yx��2~��yx��2~��x������x�      A  , ,���������������2~������2~���������      A  , ,��2~��x���2~������3(������3(��x���2~��x�      B  , ,�����{D�����{������{������{D�����{D      B  , ,�����|������}B�����}B�����|������|�      B  , ,�����}������~������~������}������}�      B  , ,�����@�����������������@�����@      B  , ,�������������>������>��������������      B  , ,�����������������������������������      B  , ,������<��������������������<������<      B  , ,�������������:������:��������������      B  , ,�����������������������������������      B  , ,������8��������������������8������8      B  , ,�������������6������6��������������      B  , ,��C��x���C��yx�����yx�����x���C��x�      B  , ,��C�����C�������������������C���      B  , ,�����x������yx��A��yx��A��x������x�      B  , ,���������������A������A���������      B  , ,�����x������yx�����yx�����x������x�      B  , ,��������������������������������      B  , ,��?��x���?��yx�����yx�����x���?��x�      B  , ,��?�����?�������������������?���      B  , ,��	���x���	���yx��
=��yx��
=��x���	���x�      B  , ,��	������	�������
=������
=�����	����      B  , ,��
���x���
���yx�����yx�����x���
���x�      B  , ,��
������
��������������������
����      B  , ,��;��x���;��yx�����yx�����x���;��x�      B  , ,��;�����;�������������������;���      B  , ,�����x������yx��9��yx��9��x������x�      B  , ,���������������9������9���������      B  , ,�����x������yx�����yx�����x������x�      B  , ,��������������������������������      B  , ,��7��x���7��yx�����yx�����x���7��x�      B  , ,��7�����7�������������������7���      B  , ,�����x������yx��5��yx��5��x������x�      B  , ,���������������5������5���������      B  , ,�����x������yx�����yx�����x������x�      B  , ,��������������������������������      B  , ,��3��x���3��yx�����yx�����x���3��x�      B  , ,��3�����3�������������������3���      B  , ,�����x������yx��1��yx��1��x������x�      B  , ,���������������1������1���������      B  , ,�����x������yx�����yx�����x������x�      B  , ,��������������������������������      B  , ,��/��x���/��yx�����yx�����x���/��x�      B  , ,��/�����/�������������������/���      B  , ,�����x������yx��-��yx��-��x������x�      B  , ,���������������-������-���������      B  , ,�����x������yx�����yx�����x������x�      B  , ,��������������������������������      B  , ,��+��x���+��yx�����yx�����x���+��x�      B  , ,��+�����+�������������������+���      B  , ,����x�����yx��)��yx��)��x�����x�      B  , ,�������������)������)��������      B  , ,�����x������yx��}��yx��}��x������x�      B  , ,���������������}������}���������      B  , ,�� '��x��� '��yx�� ���yx�� ���x��� '��x�      B  , ,�� '����� '������ ������� ������ '���      B  , ,��!{��x���!{��yx��"%��yx��"%��x���!{��x�      B  , ,��!{�����!{������"%������"%�����!{���      B  , ,��"���x���"���yx��#y��yx��#y��x���"���x�      B  , ,��"������"�������#y������#y�����"����      B  , ,��$#��x���$#��yx��$���yx��$���x���$#��x�      B  , ,��$#�����$#������$�������$������$#���      B  , ,��%w��x���%w��yx��&!��yx��&!��x���%w��x�      B  , ,��%w�����%w������&!������&!�����%w���      B  , ,��&���x���&���yx��'u��yx��'u��x���&���x�      B  , ,��&������&�������'u������'u�����&����      B  , ,��(��x���(��yx��(���yx��(���x���(��x�      B  , ,��(�����(������(�������(������(���      B  , ,��)s��x���)s��yx��*��yx��*��x���)s��x�      B  , ,��)s�����)s������*������*�����)s���      B  , ,��*���x���*���yx��+q��yx��+q��x���*���x�      B  , ,��*������*�������+q������+q�����*����      B  , ,��,��x���,��yx��,���yx��,���x���,��x�      B  , ,��,�����,������,�������,������,���      B  , ,��-o��x���-o��yx��.��yx��.��x���-o��x�      B  , ,��-o�����-o������.������.�����-o���      B  , ,��.���x���.���yx��/m��yx��/m��x���.���x�      B  , ,��.������.�������/m������/m�����.����      B  , ,��0��x���0��yx��0���yx��0���x���0��x�      B  , ,��0�����0������0�������0������0���      B  , ,��2~��{D��2~��{���3(��{���3(��{D��2~��{D      B  , ,��2~��|���2~��}B��3(��}B��3(��|���2~��|�      B  , ,��2~��}���2~��~���3(��~���3(��}���2~��}�      B  , ,��2~��@��2~�����3(�����3(��@��2~��@      B  , ,��2~������2~���>��3(���>��3(������2~����      B  , ,��2~������2~������3(������3(������2~����      B  , ,��2~���<��2~������3(������3(���<��2~���<      B  , ,��2~������2~���:��3(���:��3(������2~����      B  , ,��2~������2~������3(������3(������2~����      B  , ,��2~���8��2~������3(������3(���8��2~���8      B  , ,��2~������2~���6��3(���6��3(������2~����      B  , ,�����{������|f�����|f�����{������{�      B  , ,�����������������������������������      B  , ,��������������������������������      B  , ,��(~��{���(~��|f��0N��|f��0N��{���(~��{�      B  , ,��(~������(~������0N������0N������(~����      B  , ,��(~�����(~������0N������0N�����(~���      �   ,��1��y#��1���W��2����W��2���y#��1��y#      B   ,�����{X�����|���(j��|���(j��{X�����{X      B   ,����������������(j������(j�����������      B   ,�������������"��(j���"��(j�����������      V   ,�����y����������1f������1f��y������y�     �     0�     0 *sky130_fd_pr__res_high_po_0p35_S6WM55     B   ,��bX������bX���5��c����5��c�������bX����      B   ,��h�������h����5��i����5��i�������h�����      B   ,��n�������n����5��p"���5��p"������n�����      B   ,��t�������t����5��vX���5��vX������t�����      B   ,��{0������{0���5��|����5��|�������{0����      B   ,���f�������f���5�������5�����������f����      B   ,���������������5�������5����������������      B   ,���������������5���0���5���0������������      _   ,��a����n��a�������d������d���n��a����n      _   ,��h/���n��h/������jK������jK���n��h/���n      _   ,��ne���n��ne������p�������p����n��ne���n      _   ,��t����n��t�������v�������v����n��t����n      _   ,��z����n��z�������|�������|����n��z����n      _   ,������n����������#�������#���n������n      _   ,���=���n���=�������Y�������Y���n���=���n      _   ,���s���n���s�������������������n���s���n      C   ,��_������_����������������������_����      C   ,��_�������_������`x�����`x������_�����      C   ,��bX������bX���5��c����5��c�������bX����      C   ,��h�������h����5��i����5��i�������h�����      C   ,��n�������n����5��p"���5��p"������n�����      C   ,��t�������t����5��vX���5��vX������t�����      C   ,��{0������{0���5��|����5��|�������{0����      C   ,���f�������f���5�������5�����������f����      C   ,���������������5�������5����������������      C   ,���������������5���0���5���0������������      C   ,��bX������bX���=��c����=��c�������bX����      C   ,��h�������h����=��i����=��i�������h�����      C   ,��n�������n����=��p"���=��p"������n�����      C   ,��t�������t����=��vX���=��vX������t�����      C   ,��{0������{0���=��|����=��|�������{0����      C   ,���f�������f���=�������=�����������f����      C   ,���������������=�������=����������������      C   ,���������������=���0���=���0������������      C   ,�����������������������������������      C   ,��_����C��_��������������������C��_����C      D   ,��b�������b������c������c�������b�����      D   ,��h�������h������i������i�������h�����      D   ,��n�������n������o������o�������n�����      D   ,��u,������u,�����v&�����v&������u,����      D   ,��{b������{b�����|\�����|\������{b����      D   ,��������������������������������������      D   ,��������������������������������������      D   ,�����������������������������������      D   ,��b�������b����$��c����$��c�������b�����      D   ,��h�������h����$��i����$��i�������h�����      D   ,��n�������n����$��o����$��o�������n�����      D   ,��u,������u,���$��v&���$��v&������u,����      D   ,��{b������{b���$��|\���$��|\������{b����      D   ,���������������$�������$����������������      D   ,���������������$�������$����������������      D   ,�������������$�������$���������������      C  , ,��b����'��b�������c\������c\���'��b����'      C  , ,��h����'��h�������i�������i����'��h����'      C  , ,��o���'��o������o�������o����'��o���'      C  , ,��uT���'��uT������u�������u����'��uT���'      C  , ,��{����'��{�������|4������|4���'��{����'      C  , ,�������'�����������j�������j���'�������'      C  , ,�������'�����������������������'�������'      C  , ,���,���'���,�������������������'���,���'      C  , ,��b�������b����i��c\���i��c\������b�����      C  , ,��h�������h����i��i����i��i�������h�����      C  , ,��o������o���i��o����i��o�������o����      C  , ,��uT������uT���i��u����i��u�������uT����      C  , ,��{�������{����i��|4���i��|4������{�����      C  , ,���������������i���j���i���j������������      C  , ,���������������i�������i����������������      C  , ,���,�������,���i�������i�����������,����      C  , ,��b����W��b������c\�����c\���W��b����W      C  , ,��h����W��h������i������i����W��h����W      C  , ,��o���W��o�����o������o����W��o���W      C  , ,��uT���W��uT�����u������u����W��uT���W      C  , ,��{����W��{������|4�����|4���W��{����W      C  , ,�������W����������j������j���W�������W      C  , ,�������W���������������������W�������W      C  , ,���,���W���,�����������������W���,���W      C  , ,��b�������b������c\�����c\������b�����      C  , ,��h�������h������i������i�������h�����      C  , ,��o������o�����o������o�������o����      C  , ,��uT������uT�����u������u�������uT����      C  , ,��{�������{������|4�����|4������{�����      C  , ,������������������j������j������������      C  , ,��������������������������������������      C  , ,���,�������,���������������������,����      C  , ,��b������b����1��c\���1��c\�����b����      C  , ,��h������h����1��i����1��i������h����      C  , ,��o�����o���1��o����1��o������o���      C  , ,��uT�����uT���1��u����1��u������uT���      C  , ,��{������{����1��|4���1��|4�����{����      C  , ,��������������1���j���1���j����������      C  , ,��������������1�������1��������������      C  , ,���,������,���1�������1����������,���      C  , ,��b������b�������c\������c\�����b����      C  , ,��h������h�������i�������i������h����      C  , ,��o�����o������o�������o������o���      C  , ,��uT�����uT������u�������u������uT���      C  , ,��{������{�������|4������|4�����{����      C  , ,������������������j�������j����������      C  , ,�������������������������������������      C  , ,���,������,����������������������,���      C  , ,��b����4��b�������c\������c\���4��b����4      C  , ,��h����4��h�������i�������i����4��h����4      C  , ,��o���4��o������o�������o����4��o���4      C  , ,��uT���4��uT������u�������u����4��uT���4      C  , ,��{����4��{�������|4������|4���4��{����4      C  , ,�������4�����������j�������j���4�������4      C  , ,�������4�����������������������4�������4      C  , ,���,���4���,�������������������4���,���4      C  , ,��b�������b����v��c\���v��c\������b�����      C  , ,��h�������h����v��i����v��i�������h�����      C  , ,��o������o���v��o����v��o�������o����      C  , ,��uT������uT���v��u����v��u�������uT����      C  , ,��{�������{����v��|4���v��|4������{�����      C  , ,���������������v���j���v���j������������      C  , ,���������������v�������v����������������      C  , ,���,�������,���v�������v�����������,����      C  , ,��b����d��b������c\�����c\���d��b����d      C  , ,��h����d��h������i������i����d��h����d      C  , ,��o���d��o�����o������o����d��o���d      C  , ,��uT���d��uT�����u������u����d��uT���d      C  , ,��{����d��{������|4�����|4���d��{����d      C  , ,�������d����������j������j���d�������d      C  , ,�������d���������������������d�������d      C  , ,���,���d���,�����������������d���,���d      C  , ,��b�������b���צ��c\��צ��c\������b�����      C  , ,��h�������h���צ��i���צ��i�������h�����      C  , ,��o������o��צ��o���צ��o�������o����      C  , ,��uT������uT��צ��u���צ��u�������uT����      C  , ,��{�������{���צ��|4��צ��|4������{�����      C  , ,��������������צ���j��צ���j������������      C  , ,��������������צ������צ����������������      C  , ,���,�������,��צ������צ�����������,����      C  , ,��b���Ք��b����>��c\���>��c\��Ք��b���Ք      C  , ,��h���Ք��h����>��i����>��i���Ք��h���Ք      C  , ,��o��Ք��o���>��o����>��o���Ք��o��Ք      C  , ,��uT��Ք��uT���>��u����>��u���Ք��uT��Ք      C  , ,��{���Ք��{����>��|4���>��|4��Ք��{���Ք      C  , ,������Ք�������>���j���>���j��Ք������Ք      C  , ,������Ք�������>�������>������Ք������Ք      C  , ,���,��Ք���,���>�������>������Ք���,��Ք      C  , ,��b����,��b�������c\������c\���,��b����,      C  , ,��h����,��h�������i�������i����,��h����,      C  , ,��o���,��o������o�������o����,��o���,      C  , ,��uT���,��uT������u�������u����,��uT���,      C  , ,��{����,��{�������|4������|4���,��{����,      C  , ,�������,�����������j�������j���,�������,      C  , ,�������,�����������������������,�������,      C  , ,���,���,���,�������������������,���,���,      ^   ,��_Q������_Q���<���7���<���7������_Q����      ^   ,��_Q���j��_Q������d$������d$���j��_Q���j      ^   ,��h ���j��h ������jZ������jZ���j��h ���j      ^   ,��nV���j��nV������p�������p����j��nV���j      ^   ,��t����j��t�������v�������v����j��t����j      ^   ,��z����j��z�������|�������|����j��z����j      ^   ,�������j�����������2�������2���j�������j      ^   ,���.���j���.�������h�������h���j���.���j      ^   ,���d���j���d�������7�������7���j���d���j      ^   ,��_Q������_Q���j���7���j���7������_Q����      A  , ,��_������_����������������������_����      A  , ,��_�������_������`x�����`x������_�����      A  , ,�����������������������������������      A  , ,��_����C��_��������������������C��_����C      B  , ,��xo�����xo������y������y�����xo���      B  , ,��xo���C��xo������y������y���C��xo���C      B  , ,��{�����{������{�������{������{���      B  , ,��|k�����|k������}������}�����|k���      B  , ,��}������}�������~i������~i�����}����      B  , ,�����������������������������      B  , ,���g������g��������������������g���      B  , ,������������������e�������e����������      B  , ,����������������������������������      B  , ,���c������c��������������������c���      B  , ,������������������a�������a����������      B  , ,����������������������������������      B  , ,���_������_�������	�������	������_���      B  , ,������������������]�������]����������      B  , ,����������������������������������      B  , ,���[������[��������������������[���      B  , ,������������������Y�������Y����������      B  , ,����������������������������������      B  , ,�������������D�������D���������������      B  , ,������F����������������������F������F      B  , ,�������������������������������������      B  , ,������������H�������H�������������      B  , ,������J����������������������J������J      B  , ,�����������������������������������      B  , ,������������L�������L�������������      B  , ,������N����������������������N������N      B  , ,�����������������������������������      B  , ,������������P�������P�������������      B  , ,������R����������������������R������R      B  , ,�����������������������������������      B  , ,������������T�������T�������������      B  , ,������V������ ������� �������V������V      B  , ,��y������y�������zm������zm�����y����      B  , ,��{������{�������|>������|>�����{����      B  , ,������������������t�������t����������      B  , ,�������������������������������������      B  , ,���"������"����������������������"���      B  , ,��_����F��_�������`x������`x���F��_����F      B  , ,��d������d�������e-������e-�����d����      B  , ,��_�������_�������`x������`x������_�����      B  , ,��e������e�������f�������f������e����      B  , ,��_������_����H��`x���H��`x�����_����      B  , ,��g+�����g+������g�������g������g+���      B  , ,��_����J��_�������`x������`x���J��_����J      B  , ,��h�����h������i)������i)�����h���      B  , ,��_�������_������`x�����`x������_�����      B  , ,��i������i�������j}������j}�����i����      B  , ,��_������_����L��`x���L��`x�����_����      B  , ,��k'�����k'������k�������k������k'���      B  , ,��_����N��_�������`x������`x���N��_����N      B  , ,��l{�����l{������m%������m%�����l{���      B  , ,��_�������_������`x�����`x������_�����      B  , ,��m������m�������ny������ny�����m����      B  , ,��_������_����P��`x���P��`x�����_����      B  , ,��o#�����o#������o�������o������o#���      B  , ,��_����R��_�������`x������`x���R��_����R      B  , ,��pw�����pw������q!������q!�����pw���      B  , ,��_�������_������`x�����`x������_�����      B  , ,��q������q�������ru������ru�����q����      B  , ,��_������_����T��`x���T��`x�����_����      B  , ,��s�����s������s�������s������s���      B  , ,��_����V��_���� ��`x��� ��`x���V��_����V      B  , ,��ts�����ts������u������u�����ts���      B  , ,��u������u�������vq������vq�����u����      B  , ,��b������b�������cf������cf�����b����      B  , ,��h������h�������i�������i������h����      B  , ,��o�����o������o�������o������o���      B  , ,��uJ�����uJ������v������v�����uJ���      B  , ,��w�����w������w�������w������w���      B  , ,��a������a�������b�������b������a����      B  , ,��_�������_����D��`x���D��`x������_�����      B  , ,��c/�����c/������c�������c������c/���      B  , ,��_������_���ٸ��`x��ٸ��`x�����_����      B  , ,��_���׺��_����d��`x���d��`x��׺��_���׺      B  , ,��_����f��_������`x�����`x���f��_����f      B  , ,��_������_���ռ��`x��ռ��`x�����_����      B  , ,��_���Ӿ��_����h��`x���h��`x��Ӿ��_���Ӿ      B  , ,��a����C��a�������b�������b����C��a����C      B  , ,��c/���C��c/������c�������c����C��c/���C      B  , ,��d����C��d�������e-������e-���C��d����C      B  , ,��e����C��e�������f�������f����C��e����C      B  , ,��g+���C��g+������g�������g����C��g+���C      B  , ,��h���C��h������i)������i)���C��h���C      B  , ,��i����C��i�������j}������j}���C��i����C      B  , ,��k'���C��k'������k�������k����C��k'���C      B  , ,��l{���C��l{������m%������m%���C��l{���C      B  , ,��m����C��m�������ny������ny���C��m����C      B  , ,��o#���C��o#������o�������o����C��o#���C      B  , ,��pw���C��pw������q!������q!���C��pw���C      B  , ,��q����C��q�������ru������ru���C��q����C      B  , ,��s���C��s������s�������s����C��s���C      B  , ,��ts���C��ts������u������u���C��ts���C      B  , ,��u����C��u�������vq������vq���C��u����C      B  , ,��w���C��w������w�������w����C��w���C      B  , ,��_������_������`x�����`x�����_����      B  , ,��_������_����X��`x���X��`x�����_����      B  , ,��_����Z��_������`x�����`x���Z��_����Z      B  , ,��_������_������`x�����`x�����_����      B  , ,��_���߲��_����\��`x���\��`x��߲��_���߲      B  , ,��_����^��_������`x�����`x���^��_����^      B  , ,��_����
��_���ݴ��`x��ݴ��`x���
��_����
      B  , ,��_���۶��_����`��`x���`��`x��۶��_���۶      B  , ,��_����b��_������`x�����`x���b��_����b      B  , ,��b������b�������cf������cf�����b����      B  , ,��h������h�������i�������i������h����      B  , ,��o�����o������o�������o������o���      B  , ,��uJ�����uJ������v������v�����uJ���      B  , ,��������������������������������      B  , ,������b��������������������b������b      B  , ,��y����C��y�������zm������zm���C��y����C      B  , ,��{���C��{������{�������{����C��{���C      B  , ,��|k���C��|k������}������}���C��|k���C      B  , ,��}����C��}�������~i������~i���C��}����C      B  , ,�����C�������������������C�����C      B  , ,���g���C���g�����������������C���g���C      B  , ,�������C�����������e�������e���C�������C      B  , ,������C����������������������C������C      B  , ,���c���C���c�����������������C���c���C      B  , ,�������C�����������a�������a���C�������C      B  , ,������C����������������������C������C      B  , ,���_���C���_�������	�������	���C���_���C      B  , ,�������C�����������]�������]���C�������C      B  , ,������C����������������������C������C      B  , ,���[���C���[�����������������C���[���C      B  , ,�������C�����������Y�������Y���C�������C      B  , ,������C����������������������C������C      B  , ,�����߲������\�������\������߲�����߲      B  , ,�����������ٸ������ٸ�������������      B  , ,������Z��������������������Z������Z      B  , ,�����׺������d�������d������׺�����׺      B  , ,������^��������������������^������^      B  , ,������f��������������������f������f      B  , ,������������X�������X�������������      B  , ,�����������ռ������ռ�������������      B  , ,������
�����ݴ������ݴ�������
������
      B  , ,�����Ӿ������h�������h������Ӿ�����Ӿ      B  , ,��������������������������������      B  , ,�����۶������`�������`������۶�����۶      B  , ,��{������{�������|>������|>�����{����      B  , ,������������������t�������t����������      B  , ,�������������������������������������      B  , ,���"������"����������������������"���      �   ,��`#��ј��`#���j���e���j���e��ј��`#��ј      B   ,��bX�����bX�����c������c������bX���      B   ,��h������h������i������i������h����      B   ,��n������n������p"�����p"�����n����      B   ,��t������t������vX�����vX�����t����      B   ,��{0�����{0�����|������|������{0���      B   ,���f������f��������������������f���      B   ,�����������������������������������      B   ,�����������������0������0����������      V   ,��`������`����������������������`����     �     0�     0 *sky130_fd_pr__res_high_po_0p35_5T4P9C     B   ,���������������J���M���J���M������������      B   ,��%������%���J������J���������%����      B   ,��
[������
[���J������J���������
[����      B   ,�������������J������J��������������      B   ,�������������J��%���J��%�����������      B   ,�������������J��[���J��[�����������      B   ,��#3������#3���J��$����J��$�������#3����      B   ,��)i������)i���J��*����J��*�������)i����      _   ,�������k�����������������������k�������k      _   ,������k��������������������k������k      _   ,��	����k��	����������������k��	����k      _   ,��2���k��2������N������N���k��2���k      _   ,��h���k��h�����������������k��h���k      _   ,������k��������������������k������k      _   ,��"����k��"�������$�������$����k��"����k      _   ,��)
���k��)
������+&������+&���k��)
���k      C   ,���e���*���e������-Q������-Q���*���e���*      C   ,���e�������e���*������*����������e����      C   ,���������������J���M���J���M������������      C   ,��%������%���J������J���������%����      C   ,��
[������
[���J������J���������
[����      C   ,�������������J������J��������������      C   ,�������������J��%���J��%�����������      C   ,�������������J��[���J��[�����������      C   ,��#3������#3���J��$����J��$�������#3����      C   ,��)i������)i���J��*����J��*�������)i����      C   ,���������������:���M���:���M������������      C   ,��%������%���:������:���������%����      C   ,��
[������
[���:������:���������
[����      C   ,�������������:������:��������������      C   ,�������������:��%���:��%�����������      C   ,�������������:��[���:��[�����������      C   ,��#3������#3���:��$����:��$�������#3����      C   ,��)i������)i���:��*����:��*�������)i����      C   ,��,�������,����*��-Q���*��-Q������,�����      C   ,���e���@���e������-Q������-Q���@���e���@      D   ,���!�������!���,������,����������!����      D   ,��W������W���,��Q���,��Q������W����      D   ,��
�������
����,������,���������
�����      D   ,�������������,������,��������������      D   ,�������������,������,��������������      D   ,��/������/���,��)���,��)������/����      D   ,��#e������#e���,��$_���,��$_������#e����      D   ,��)�������)����,��*����,��*�������)�����      D   ,���!�������!���!������!����������!����      D   ,��W������W���!��Q���!��Q������W����      D   ,��
�������
����!������!���������
�����      D   ,�������������!������!��������������      D   ,�������������!������!��������������      D   ,��/������/���!��)���!��)������/����      D   ,��#e������#e���!��$_���!��$_������#e����      D   ,��)�������)����!��*����!��*�������)�����      C  , ,���I���<���I�������������������<���I���<      C  , ,�����<��������)������)���<�����<      C  , ,��
����<��
�������_������_���<��
����<      C  , ,������<��������������������<������<      C  , ,��!���<��!�����������������<��!���<      C  , ,��W���<��W���������������<��W���<      C  , ,��#����<��#�������$7������$7���<��#����<      C  , ,��)����<��)�������*m������*m���<��)����<      C  , ,���I�������I���~�������~�����������I����      C  , ,�����������~��)���~��)����������      C  , ,��
�������
����~��_���~��_������
�����      C  , ,�������������~������~��������������      C  , ,��!������!���~������~���������!����      C  , ,��W������W���~�����~��������W����      C  , ,��#�������#����~��$7���~��$7������#�����      C  , ,��)�������)����~��*m���~��*m������)�����      C  , ,���I���l���I�����������������l���I���l      C  , ,�����l�������)�����)���l�����l      C  , ,��
����l��
������_�����_���l��
����l      C  , ,������l������������������l������l      C  , ,��!���l��!���������������l��!���l      C  , ,��W���l��W�������������l��W���l      C  , ,��#����l��#������$7�����$7���l��#����l      C  , ,��)����l��)������*m�����*m���l��)����l      C  , ,���I������I��������������������I���      C  , ,������������)�����)��������      C  , ,��
������
������_�����_�����
����      C  , ,������������������������������      C  , ,��!�����!�����������������!���      C  , ,��W�����W���������������W���      C  , ,��#������#������$7�����$7�����#����      C  , ,��)������)������*m�����*m�����)����      C  , ,���I������I���F�������F����������I���      C  , ,����������F��)���F��)��������      C  , ,��
������
����F��_���F��_�����
����      C  , ,������������F������F������������      C  , ,��!�����!���F������F��������!���      C  , ,��W�����W���F�����F�������W���      C  , ,��#������#����F��$7���F��$7�����#����      C  , ,��)������)����F��*m���F��*m�����)����      C  , ,���I���4���I�������������������4���I���4      C  , ,�����4��������)������)���4�����4      C  , ,��
����4��
�������_������_���4��
����4      C  , ,������4��������������������4������4      C  , ,��!���4��!�����������������4��!���4      C  , ,��W���4��W���������������4��W���4      C  , ,��#����4��#�������$7������$7���4��#����4      C  , ,��)����4��)�������*m������*m���4��)����4      C  , ,���I���1���I�������������������1���I���1      C  , ,�����1��������)������)���1�����1      C  , ,��
����1��
�������_������_���1��
����1      C  , ,������1��������������������1������1      C  , ,��!���1��!�����������������1��!���1      C  , ,��W���1��W���������������1��W���1      C  , ,��#����1��#�������$7������$7���1��#����1      C  , ,��)����1��)�������*m������*m���1��)����1      C  , ,���I�������I���s�������s�����������I����      C  , ,�����������s��)���s��)����������      C  , ,��
�������
����s��_���s��_������
�����      C  , ,�������������s������s��������������      C  , ,��!������!���s������s���������!����      C  , ,��W������W���s�����s��������W����      C  , ,��#�������#����s��$7���s��$7������#�����      C  , ,��)�������)����s��*m���s��*m������)�����      C  , ,���I���a���I�����������������a���I���a      C  , ,�����a�������)�����)���a�����a      C  , ,��
����a��
������_�����_���a��
����a      C  , ,������a������������������a������a      C  , ,��!���a��!���������������a��!���a      C  , ,��W���a��W�������������a��W���a      C  , ,��#����a��#������$7�����$7���a��#����a      C  , ,��)����a��)������*m�����*m���a��)����a      C  , ,���I�������I��ڣ������ڣ�����������I����      C  , ,����������ڣ��)��ڣ��)����������      C  , ,��
�������
���ڣ��_��ڣ��_������
�����      C  , ,������������ڣ�����ڣ��������������      C  , ,��!������!��ڣ�����ڣ���������!����      C  , ,��W������W��ڣ����ڣ��������W����      C  , ,��#�������#���ڣ��$7��ڣ��$7������#�����      C  , ,��)�������)���ڣ��*m��ڣ��*m������)�����      C  , ,���I��ؑ���I���;�������;������ؑ���I��ؑ      C  , ,����ؑ�����;��)���;��)��ؑ����ؑ      C  , ,��
���ؑ��
����;��_���;��_��ؑ��
���ؑ      C  , ,�����ؑ������;������;�����ؑ�����ؑ      C  , ,��!��ؑ��!���;������;�����ؑ��!��ؑ      C  , ,��W��ؑ��W���;�����;����ؑ��W��ؑ      C  , ,��#���ؑ��#����;��$7���;��$7��ؑ��#���ؑ      C  , ,��)���ؑ��)����;��*m���;��*m��ؑ��)���ؑ      C  , ,���I���)���I�������������������)���I���)      C  , ,�����)��������)������)���)�����)      C  , ,��
����)��
�������_������_���)��
����)      C  , ,������)��������������������)������)      C  , ,��!���)��!�����������������)��!���)      C  , ,��W���)��W���������������)��W���)      C  , ,��#����)��#�������$7������$7���)��#����)      C  , ,��)����)��)�������*m������*m���)��)����)      ^   ,���������������Q��-����Q��-�������������      ^   ,�������g�����������������������g�������g      ^   ,������g��������������������g������g      ^   ,��	����g��	�������'������'���g��	����g      ^   ,��#���g��#������]������]���g��#���g      ^   ,��Y���g��Y�����������������g��Y���g      ^   ,������g��������������������g������g      ^   ,��"����g��"�������$�������$����g��"����g      ^   ,��(����g��(�������-�������-����g��(����g      ^   ,���������������g��-����g��-�������������      A  , ,���e���*���e������-Q������-Q���*���e���*      A  , ,���e�������e���*������*����������e����      A  , ,��,�������,����*��-Q���*��-Q������,�����      A  , ,���e���@���e������-Q������-Q���@���e���@      B  , ,�����*�������������������*�����*      B  , ,���e������e���_������_���������e���      B  , ,��,������,����_��-Q���_��-Q�����,����      B  , ,�����@�������������������@�����@      B  , ,��V���*��V������ ������ ���*��V���*      B  , ,������*���������T������T���*������*      B  , ,������*��������������������*������*      B  , ,��R���*��R�����������������*��R���*      B  , ,������*���������P������P���*������*      B  , ,������*��������� ������� ����*������*      B  , ,��!N���*��!N������!�������!����*��!N���*      B  , ,��"����*��"�������#L������#L���*��"����*      B  , ,��#����*��#�������$�������$����*��#����*      B  , ,��%J���*��%J������%�������%����*��%J���*      B  , ,��&����*��&�������'H������'H���*��&����*      B  , ,��'����*��'�������(�������(����*��'����*      B  , ,��)F���*��)F������)�������)����*��)F���*      B  , ,��*����*��*�������+D������+D���*��*����*      B  , ,��,�������,����O��-Q���O��-Q������,�����      B  , ,��,����Q��,�������-Q������-Q���Q��,����Q      B  , ,��,�������,�������-Q������-Q������,�����      B  , ,��,������,����S��-Q���S��-Q�����,����      B  , ,��,����U��,�������-Q������-Q���U��,����U      B  , ,��,������,������-Q�����-Q�����,����      B  , ,��,������,����W��-Q���W��-Q�����,����      B  , ,��,����Y��,������-Q�����-Q���Y��,����Y      B  , ,��,������,������-Q�����-Q�����,����      B  , ,��,������,����[��-Q���[��-Q�����,����      B  , ,��,����]��,������-Q�����-Q���]��,����]      B  , ,��,����	��,������-Q�����-Q���	��,����	      B  , ,��Z���*��Z���������������*��Z���*      B  , ,������*���������X������X���*������*      B  , ,�����*�������������������*�����*      B  , ,�����*�������������������*�����*      B  , ,��M���*��M���������������*��M���*      B  , ,��#����*��#�������$A������$A���*��#����*      B  , ,��)����*��)�������*w������*w���*��)����*      B  , ,���e���Q���e�����������������Q���e���Q      B  , ,�� ���*�� ������ ������� ����*�� ���*      B  , ,���e�������e���������������������e����      B  , ,��n���*��n���������������*��n���*      B  , ,���e������e���S������S���������e���      B  , ,������*���������l������l���*������*      B  , ,���e���U���e�����������������U���e���U      B  , ,�����*�������������������*�����*      B  , ,���e������e������������������e���      B  , ,��j���*��j���������������*��j���*      B  , ,���e������e���W������W���������e���      B  , ,������*���������h������h���*������*      B  , ,���e���Y���e���������������Y���e���Y      B  , ,�����*�������������������*�����*      B  , ,���e������e������������������e���      B  , ,��	f���*��	f������
������
���*��	f���*      B  , ,���e������e���[������[���������e���      B  , ,��
����*��
�������d������d���*��
����*      B  , ,���e���]���e���������������]���e���]      B  , ,�����*�������������������*�����*      B  , ,���e���	���e���������������	���e���	      B  , ,��b���*��b���������������*��b���*      B  , ,������*���������`������`���*������*      B  , ,��
���*��
�����������������*��
���*      B  , ,��^���*��^���������������*��^���*      B  , ,���?���*���?�������������������*���?���*      B  , ,��u���*��u������3������3���*��u���*      B  , ,��
����*��
�������i������i���*��
����*      B  , ,������*��������������������*������*      B  , ,������*���������\������\���*������*      B  , ,���r���*���r�����������������*���r���*      B  , ,���e�������e���O������O����������e����      B  , ,�������*�����������p�������p���*�������*      B  , ,���e���m���e���������������m���e���m      B  , ,���e������e��������������������e���      B  , ,���e�������e���o������o����������e����      B  , ,���r���@���r�����������������@���r���@      B  , ,�������@�����������p�������p���@�������@      B  , ,�� ���@�� ������ ������� ����@�� ���@      B  , ,��n���@��n���������������@��n���@      B  , ,������@���������l������l���@������@      B  , ,�����@�������������������@�����@      B  , ,��j���@��j���������������@��j���@      B  , ,������@���������h������h���@������@      B  , ,�����@�������������������@�����@      B  , ,��	f���@��	f������
������
���@��	f���@      B  , ,��
����@��
�������d������d���@��
����@      B  , ,�����@�������������������@�����@      B  , ,��b���@��b���������������@��b���@      B  , ,������@���������`������`���@������@      B  , ,��
���@��
�����������������@��
���@      B  , ,��^���@��^���������������@��^���@      B  , ,������@���������\������\���@������@      B  , ,���e���a���e���������������a���e���a      B  , ,���e������e������������������e���      B  , ,���e������e���c������c���������e���      B  , ,���e���e���e���������������e���e���e      B  , ,���e������e������������������e���      B  , ,���e��޽���e���g������g�����޽���e��޽      B  , ,���e���i���e���������������i���e���i      B  , ,���e������e��ܿ�����ܿ���������e���      B  , ,���e�������e���k������k����������e����      B  , ,���?������?����������������������?���      B  , ,��u�����u������3������3�����u���      B  , ,��
������
�������i������i�����
����      B  , ,��������������������������������      B  , ,��Z���@��Z���������������@��Z���@      B  , ,������@���������X������X���@������@      B  , ,�����@�������������������@�����@      B  , ,��V���@��V������ ������ ���@��V���@      B  , ,������@���������T������T���@������@      B  , ,������@��������������������@������@      B  , ,��R���@��R�����������������@��R���@      B  , ,������@���������P������P���@������@      B  , ,������@��������� ������� ����@������@      B  , ,��!N���@��!N������!�������!����@��!N���@      B  , ,��"����@��"�������#L������#L���@��"����@      B  , ,��#����@��#�������$�������$����@��#����@      B  , ,��%J���@��%J������%�������%����@��%J���@      B  , ,��&����@��&�������'H������'H���@��&����@      B  , ,��'����@��'�������(�������(����@��'����@      B  , ,��)F���@��)F������)�������)����@��)F���@      B  , ,��*����@��*�������+D������+D���@��*����@      B  , ,��,������,������-Q�����-Q�����,����      B  , ,��,����m��,������-Q�����-Q���m��,����m      B  , ,��,������,����c��-Q���c��-Q�����,����      B  , ,��,������,�������-Q������-Q�����,����      B  , ,��,���޽��,����g��-Q���g��-Q��޽��,���޽      B  , ,��,�������,����o��-Q���o��-Q������,�����      B  , ,��,������,������-Q�����-Q�����,����      B  , ,��,����i��,������-Q�����-Q���i��,����i      B  , ,��,����e��,������-Q�����-Q���e��,����e      B  , ,��,������,���ܿ��-Q��ܿ��-Q�����,����      B  , ,��,����a��,������-Q�����-Q���a��,����a      B  , ,��,�������,����k��-Q���k��-Q������,�����      B  , ,�����������������������������      B  , ,��M�����M�����������������M���      B  , ,��#������#�������$A������$A�����#����      B  , ,��)������)�������*w������*w�����)����      �   ,������ԕ���������,������,���ԕ������ԕ      B   ,������������������M������M������������      B   ,��%������%������������������%����      B   ,��
[������
[������������������
[����      B   ,���������������������������������      B   ,���������������%�����%�����������      B   ,���������������[�����[�����������      B   ,��#3������#3�����$������$�������#3����      B   ,��)i������)i�����*������*�������)i����      V   ,���#������#�����,������,�������#���     �     0�     0 *sky130_fd_pr__res_xhigh_po_0p35_Y3K8LK    B   ,��I�  I��I�  "���J�  "���J�  I��I�  I      B   ,��O�  I��O�  "���Q  "���Q  I��O�  I      B   ,��U�  I��U�  "���WJ  "���WJ  I��U�  I      B   ,��\"  I��\"  "���]�  "���]�  I��\"  I      B   ,��bX  I��bX  "���c�  "���c�  I��bX  I      B   ,��h�  I��h�  "���i�  "���i�  I��h�  I      _   ,��I!  ���I!  #(��K=  #(��K=  ���I!  �      _   ,��OW  ���OW  #(��Qs  #(��Qs  ���OW  �      _   ,��U�  ���U�  #(��W�  #(��W�  ���U�  �      _   ,��[�  ���[�  #(��]�  #(��]�  ���[�  �      _   ,��a�  ���a�  #(��d  #(��d  ���a�  �      _   ,��h/  ���h/  #(��jK  #(��jK  ���h/  �      C   ,��F�  $���F�  %S��lv  %S��lv  $���F�  $�      C   ,��F�   i��F�  $���G�  $���G�   i��F�   i      C   ,��I�  Y��I�  "���J�  "���J�  Y��I�  Y      C   ,��O�  Y��O�  "���Q  "���Q  Y��O�  Y      C   ,��U�  Y��U�  "���WJ  "���WJ  Y��U�  Y      C   ,��\"  Y��\"  "���]�  "���]�  Y��\"  Y      C   ,��bX  Y��bX  "���c�  "���c�  Y��bX  Y      C   ,��h�  Y��h�  "���i�  "���i�  Y��h�  Y      C   ,��I�  I��I�  
���J�  
���J�  I��I�  I      C   ,��O�  I��O�  
���Q  
���Q  I��O�  I      C   ,��U�  I��U�  
���WJ  
���WJ  I��U�  I      C   ,��\"  I��\"  
���]�  
���]�  I��\"  I      C   ,��bX  I��bX  
���c�  
���c�  I��bX  I      C   ,��h�  I��h�  
���i�  
���i�  I��h�  I      C   ,��k�   i��k�  $���lv  $���lv   i��k�   i      C   ,��F�������F�   i��lv   i��lv������F�����      D   ,��I�  r��I�  "���J�  "���J�  r��I�  r      D   ,��O�  r��O�  "���P�  "���P�  r��O�  r      D   ,��V  r��V  "���W  "���W  r��V  r      D   ,��\T  r��\T  "���]N  "���]N  r��\T  r      D   ,��b�  r��b�  "���c�  "���c�  r��b�  r      D   ,��h�  r��h�  "���i�  "���i�  r��h�  r      D   ,��I�  g��I�  
���J�  
���J�  g��I�  g      D   ,��O�  g��O�  
���P�  
���P�  g��O�  g      D   ,��V  g��V  
���W  
���W  g��V  g      D   ,��\T  g��\T  
���]N  
���]N  g��\T  g      D   ,��b�  g��b�  
���c�  
���c�  g��b�  g      D   ,��h�  g��h�  
���i�  
���i�  g��h�  g      C  , ,��I�  !���I�  "e��J�  "e��J�  !���I�  !�      C  , ,��P  !���P  "e��P�  "e��P�  !���P  !�      C  , ,��VF  !���VF  "e��V�  "e��V�  !���VF  !�      C  , ,��\|  !���\|  "e��]&  "e��]&  !���\|  !�      C  , ,��b�  !���b�  "e��c\  "e��c\  !���b�  !�      C  , ,��h�  !���h�  "e��i�  "e��i�  !���h�  !�      C  , ,��I�   S��I�   ���J�   ���J�   S��I�   S      C  , ,��P   S��P   ���P�   ���P�   S��P   S      C  , ,��VF   S��VF   ���V�   ���V�   S��VF   S      C  , ,��\|   S��\|   ���]&   ���]&   S��\|   S      C  , ,��b�   S��b�   ���c\   ���c\   S��b�   S      C  , ,��h�   S��h�   ���i�   ���i�   S��h�   S      C  , ,��I�  ���I�  ���J�  ���J�  ���I�  �      C  , ,��P  ���P  ���P�  ���P�  ���P  �      C  , ,��VF  ���VF  ���V�  ���V�  ���VF  �      C  , ,��\|  ���\|  ���]&  ���]&  ���\|  �      C  , ,��b�  ���b�  ���c\  ���c\  ���b�  �      C  , ,��h�  ���h�  ���i�  ���i�  ���h�  �      C  , ,��I�  ���I�  -��J�  -��J�  ���I�  �      C  , ,��P  ���P  -��P�  -��P�  ���P  �      C  , ,��VF  ���VF  -��V�  -��V�  ���VF  �      C  , ,��\|  ���\|  -��]&  -��]&  ���\|  �      C  , ,��b�  ���b�  -��c\  -��c\  ���b�  �      C  , ,��h�  ���h�  -��i�  -��i�  ���h�  �      C  , ,��I�  ��I�  ���J�  ���J�  ��I�        C  , ,��P  ��P  ���P�  ���P�  ��P        C  , ,��VF  ��VF  ���V�  ���V�  ��VF        C  , ,��\|  ��\|  ���]&  ���]&  ��\|        C  , ,��b�  ��b�  ���c\  ���c\  ��b�        C  , ,��h�  ��h�  ���i�  ���i�  ��h�        C  , ,��I�  ���I�  ]��J�  ]��J�  ���I�  �      C  , ,��P  ���P  ]��P�  ]��P�  ���P  �      C  , ,��VF  ���VF  ]��V�  ]��V�  ���VF  �      C  , ,��\|  ���\|  ]��]&  ]��]&  ���\|  �      C  , ,��b�  ���b�  ]��c\  ]��c\  ���b�  �      C  , ,��h�  ���h�  ]��i�  ]��i�  ���h�  �      C  , ,��I�  	���I�  
Z��J�  
Z��J�  	���I�  	�      C  , ,��P  	���P  
Z��P�  
Z��P�  	���P  	�      C  , ,��VF  	���VF  
Z��V�  
Z��V�  	���VF  	�      C  , ,��\|  	���\|  
Z��]&  
Z��]&  	���\|  	�      C  , ,��b�  	���b�  
Z��c\  
Z��c\  	���b�  	�      C  , ,��h�  	���h�  
Z��i�  
Z��i�  	���h�  	�      C  , ,��I�  H��I�  ���J�  ���J�  H��I�  H      C  , ,��P  H��P  ���P�  ���P�  H��P  H      C  , ,��VF  H��VF  ���V�  ���V�  H��VF  H      C  , ,��\|  H��\|  ���]&  ���]&  H��\|  H      C  , ,��b�  H��b�  ���c\  ���c\  H��b�  H      C  , ,��h�  H��h�  ���i�  ���i�  H��h�  H      C  , ,��I�  ���I�  ���J�  ���J�  ���I�  �      C  , ,��P  ���P  ���P�  ���P�  ���P  �      C  , ,��VF  ���VF  ���V�  ���V�  ���VF  �      C  , ,��\|  ���\|  ���]&  ���]&  ���\|  �      C  , ,��b�  ���b�  ���c\  ���c\  ���b�  �      C  , ,��h�  ���h�  ���i�  ���i�  ���h�  �      C  , ,��I�  x��I�  "��J�  "��J�  x��I�  x      C  , ,��P  x��P  "��P�  "��P�  x��P  x      C  , ,��VF  x��VF  "��V�  "��V�  x��VF  x      C  , ,��\|  x��\|  "��]&  "��]&  x��\|  x      C  , ,��b�  x��b�  "��c\  "��c\  x��b�  x      C  , ,��h�  x��h�  "��i�  "��i�  x��h�  x      C  , ,��I�  ��I�  ���J�  ���J�  ��I�        C  , ,��P  ��P  ���P�  ���P�  ��P        C  , ,��VF  ��VF  ���V�  ���V�  ��VF        C  , ,��\|  ��\|  ���]&  ���]&  ��\|        C  , ,��b�  ��b�  ���c\  ���c\  ��b�        C  , ,��h�  ��h�  ���i�  ���i�  ��h�        C  , ,��I�  ���I�  R��J�  R��J�  ���I�  �      C  , ,��P  ���P  R��P�  R��P�  ���P  �      C  , ,��VF  ���VF  R��V�  R��V�  ���VF  �      C  , ,��\|  ���\|  R��]&  R��]&  ���\|  �      C  , ,��b�  ���b�  R��c\  R��c\  ���b�  �      C  , ,��h�  ���h�  R��i�  R��i�  ���h�  �      ^   ,��Fy  $,��Fy  %���l�  %���l�  $,��Fy  $,      ^   ,��Fy   ���Fy  $,��KL  $,��KL   ���Fy   �      ^   ,��OH   ���OH  $,��Q�  $,��Q�   ���OH   �      ^   ,��U~   ���U~  $,��W�  $,��W�   ���U~   �      ^   ,��[�   ���[�  $,��]�  $,��]�   ���[�   �      ^   ,��a�   ���a�  $,��d$  $,��d$   ���a�   �      ^   ,��h    ���h   $,��l�  $,��l�   ���h    �      ^   ,��Fy���B��Fy   ���l�   ���l����B��Fy���B      A  , ,��F�  $���F�  %S��lv  %S��lv  $���F�  $�      A  , ,��F�   i��F�  $���G�  $���G�   i��F�   i      A  , ,��k�   i��k�  $���lv  $���lv   i��k�   i      A  , ,��F�������F�   i��lv   i��lv������F�����      B  , ,��Ya  $���Ya  %S��Z  %S��Z  $���Ya  $�      B  , ,��F�  4��F�  ���G�  ���G�  4��F�  4      B  , ,��k�  4��k�  ���lv  ���lv  4��k�  4      B  , ,��Ya������Ya   i��Z   i��Z������Ya����      B  , ,��^�  $���^�  %S��_[  %S��_[  $���^�  $�      B  , ,��`  $���`  %S��`�  %S��`�  $���`  $�      B  , ,��aY  $���aY  %S��b  %S��b  $���aY  $�      B  , ,��b�  $���b�  %S��cW  %S��cW  $���b�  $�      B  , ,��d  $���d  %S��d�  %S��d�  $���d  $�      B  , ,��eU  $���eU  %S��e�  %S��e�  $���eU  $�      B  , ,��f�  $���f�  %S��gS  %S��gS  $���f�  $�      B  , ,��g�  $���g�  %S��h�  %S��h�  $���g�  $�      B  , ,��iQ  $���iQ  %S��i�  %S��i�  $���iQ  $�      B  , ,��k�  "$��k�  "���lv  "���lv  "$��k�  "$      B  , ,��k�   ���k�  !z��lv  !z��lv   ���k�   �      B  , ,��k�  |��k�   &��lv   &��lv  |��k�  |      B  , ,��k�  (��k�  ���lv  ���lv  (��k�  (      B  , ,��k�  ���k�  ~��lv  ~��lv  ���k�  �      B  , ,��k�  ���k�  *��lv  *��lv  ���k�  �      B  , ,��k�  ,��k�  ���lv  ���lv  ,��k�  ,      B  , ,��k�  ���k�  ���lv  ���lv  ���k�  �      B  , ,��k�  ���k�  .��lv  .��lv  ���k�  �      B  , ,��k�  0��k�  ���lv  ���lv  0��k�  0      B  , ,��k�  ���k�  ���lv  ���lv  ���k�  �      B  , ,��k�  ���k�  2��lv  2��lv  ���k�  �      B  , ,��Z�  $���Z�  %S��[_  %S��[_  $���Z�  $�      B  , ,��\	  $���\	  %S��\�  %S��\�  $���\	  $�      B  , ,��]]  $���]]  %S��^  %S��^  $���]]  $�      B  , ,��\r  ���\r  "y��]0  "y��]0  ���\r  �      B  , ,��b�  ���b�  "y��cf  "y��cf  ���b�  �      B  , ,��h�  ���h�  "y��i�  "y��i�  ���h�  �      B  , ,��F�  (��F�  ���G�  ���G�  (��F�  (      B  , ,��N�  $���N�  %S��Ok  %S��Ok  $���N�  $�      B  , ,��F�  ���F�  ~��G�  ~��G�  ���F�  �      B  , ,��P  $���P  %S��P�  %S��P�  $���P  $�      B  , ,��F�  ���F�  *��G�  *��G�  ���F�  �      B  , ,��Qi  $���Qi  %S��R  %S��R  $���Qi  $�      B  , ,��F�  ,��F�  ���G�  ���G�  ,��F�  ,      B  , ,��R�  $���R�  %S��Sg  %S��Sg  $���R�  $�      B  , ,��F�  ���F�  ���G�  ���G�  ���F�  �      B  , ,��T  $���T  %S��T�  %S��T�  $���T  $�      B  , ,��F�  ���F�  .��G�  .��G�  ���F�  �      B  , ,��Ue  $���Ue  %S��V  %S��V  $���Ue  $�      B  , ,��F�  0��F�  ���G�  ���G�  0��F�  0      B  , ,��V�  $���V�  %S��Wc  %S��Wc  $���V�  $�      B  , ,��F�  ���F�  ���G�  ���G�  ���F�  �      B  , ,��X  $���X  %S��X�  %S��X�  $���X  $�      B  , ,��F�  ���F�  2��G�  2��G�  ���F�  �      B  , ,��Iq  $���Iq  %S��J  %S��J  $���Iq  $�      B  , ,��F�  "$��F�  "���G�  "���G�  "$��F�  "$      B  , ,��J�  $���J�  %S��Ko  %S��Ko  $���J�  $�      B  , ,��F�   ���F�  !z��G�  !z��G�   ���F�   �      B  , ,��I�  ���I�  "y��J�  "y��J�  ���I�  �      B  , ,��P  ���P  "y��P�  "y��P�  ���P  �      B  , ,��V<  ���V<  "y��V�  "y��V�  ���V<  �      B  , ,��L  $���L  %S��L�  %S��L�  $���L  $�      B  , ,��F�  |��F�   &��G�   &��G�  |��F�  |      B  , ,��Mm  $���Mm  %S��N  %S��N  $���Mm  $�      B  , ,��F�  ���F�  >��G�  >��G�  ���F�  �      B  , ,��F�  @��F�  ���G�  ���G�  @��F�  @      B  , ,��F�  ���F�  ���G�  ���G�  ���F�  �      B  , ,��F�  ���F�  B��G�  B��G�  ���F�  �      B  , ,��F�  D��F�  ���G�  ���G�  D��F�  D      B  , ,��Iq������Iq   i��J   i��J������Iq����      B  , ,��J�������J�   i��Ko   i��Ko������J�����      B  , ,��L������L   i��L�   i��L�������L����      B  , ,��Mm������Mm   i��N   i��N������Mm����      B  , ,��N�������N�   i��Ok   i��Ok������N�����      B  , ,��P������P   i��P�   i��P�������P����      B  , ,��Qi������Qi   i��R   i��R������Qi����      B  , ,��R�������R�   i��Sg   i��Sg������R�����      B  , ,��T������T   i��T�   i��T�������T����      B  , ,��Ue������Ue   i��V   i��V������Ue����      B  , ,��V�������V�   i��Wc   i��Wc������V�����      B  , ,��X������X   i��X�   i��X�������X����      B  , ,��F�  ���F�  ���G�  ���G�  ���F�  �      B  , ,��F�  ���F�  6��G�  6��G�  ���F�  �      B  , ,��F�  8��F�  ���G�  ���G�  8��F�  8      B  , ,��F�  ���F�  ���G�  ���G�  ���F�  �      B  , ,��F�  ���F�  :��G�  :��G�  ���F�  �      B  , ,��F�  
<��F�  
���G�  
���G�  
<��F�  
<      B  , ,��F�  ���F�  	���G�  	���G�  ���F�  �      B  , ,��I�  ���I�  
i��J�  
i��J�  ���I�  �      B  , ,��P  ���P  
i��P�  
i��P�  ���P  �      B  , ,��V<  ���V<  
i��V�  
i��V�  ���V<  �      B  , ,��k�  
<��k�  
���lv  
���lv  
<��k�  
<      B  , ,��k�  D��k�  ���lv  ���lv  D��k�  D      B  , ,��k�  ���k�  6��lv  6��lv  ���k�  �      B  , ,��Z�������Z�   i��[_   i��[_������Z�����      B  , ,��\	������\	   i��\�   i��\�������\	����      B  , ,��]]������]]   i��^   i��^������]]����      B  , ,��^�������^�   i��_[   i��_[������^�����      B  , ,��`������`   i��`�   i��`�������`����      B  , ,��aY������aY   i��b   i��b������aY����      B  , ,��b�������b�   i��cW   i��cW������b�����      B  , ,��d������d   i��d�   i��d�������d����      B  , ,��eU������eU   i��e�   i��e�������eU����      B  , ,��f�������f�   i��gS   i��gS������f�����      B  , ,��g�������g�   i��h�   i��h�������g�����      B  , ,��iQ������iQ   i��i�   i��i�������iQ����      B  , ,��k�  ���k�  	���lv  	���lv  ���k�  �      B  , ,��k�  ���k�  ���lv  ���lv  ���k�  �      B  , ,��k�  ���k�  >��lv  >��lv  ���k�  �      B  , ,��k�  ���k�  ���lv  ���lv  ���k�  �      B  , ,��k�  @��k�  ���lv  ���lv  @��k�  @      B  , ,��k�  ���k�  :��lv  :��lv  ���k�  �      B  , ,��k�  ���k�  ���lv  ���lv  ���k�  �      B  , ,��k�  8��k�  ���lv  ���lv  8��k�  8      B  , ,��k�  ���k�  B��lv  B��lv  ���k�  �      B  , ,��\r  ���\r  
i��]0  
i��]0  ���\r  �      B  , ,��b�  ���b�  
i��cf  
i��cf  ���b�  �      B  , ,��h�  ���h�  
i��i�  
i��i�  ���h�  �      �   ,��GK   ��GK  $���l!  $���l!   ��GK         B   ,��I�  
}��I�  ���J�  ���J�  
}��I�  
}      B   ,��O�  
}��O�  ���Q  ���Q  
}��O�  
}      B   ,��U�  
}��U�  ���WJ  ���WJ  
}��U�  
}      B   ,��\"  
}��\"  ���]�  ���]�  
}��\"  
}      B   ,��bX  
}��bX  ���c�  ���c�  
}��bX  
}      B   ,��h�  
}��h�  ���i�  ���i�  
}��h�  
}      O   ,��G�  ���G�  #���k�  #���k�  ���G�  �     �     0�     0 via_new$3  	   D   !     �           �       	   E   !     �           �       	   F   !     �           �       	   G   !     �           �          D  , ,   }����   }����  ����  ����   }����      D  , ,  �����  �����  S����  S����  �����      D  , ,  �����  �����  �����  �����  �����      D  , ,  =����  =����  �����  �����  =����      D  , ,  }����  }����  ����  ����  }����      D  , ,  �����  �����  S����  S����  �����      D  , ,   }���5   }����  ����  ���5   }���5      D  , ,  ����5  �����  S����  S���5  ����5      D  , ,  ����5  �����  �����  ����5  ����5      D  , ,  =���5  =����  �����  ����5  =���5      D  , ,  }���5  }����  ����  ���5  }���5      D  , ,  ����5  �����  S����  S���5  ����5      D  , ,   }���u   }���  ���  ���u   }���u      D  , ,  ����u  ����  S���  S���u  ����u      D  , ,  ����u  ����  ����  ����u  ����u      D  , ,  =���u  =���  ����  ����u  =���u      D  , ,  }���u  }���  ���  ���u  }���u      D  , ,  ����u  ����  S���  S���u  ����u      D  , ,   }����   }���K  ���K  ����   }����      D  , ,  �����  ����K  S���K  S����  �����      D  , ,  �����  ����K  ����K  �����  �����      D  , ,  =����  =���K  ����K  �����  =����      D  , ,  }����  }���K  ���K  ����  }����      D  , ,  �����  ����K  S���K  S����  �����      D  , ,   }����   }����  ����  ����   }����      D  , ,  �����  �����  S����  S����  �����      D  , ,  �����  �����  �����  �����  �����      D  , ,  =����  =����  �����  �����  =����      D  , ,  }����  }����  ����  ����  }����      D  , ,  �����  �����  S����  S����  �����      D  , ,   }���5   }����  ����  ���5   }���5      D  , ,  ����5  �����  S����  S���5  ����5      D  , ,  ����5  �����  �����  ����5  ����5      D  , ,  =���5  =����  �����  ����5  =���5      D  , ,  }���5  }����  ����  ���5  }���5      D  , ,  ����5  �����  S����  S���5  ����5      D  , ,   }���u   }���  ���  ���u   }���u      D  , ,  ����u  ����  S���  S���u  ����u      D  , ,  ����u  ����  ����  ����u  ����u      D  , ,  =���u  =���  ����  ����u  =���u      D  , ,  }���u  }���  ���  ���u  }���u      D  , ,  ����u  ����  S���  S���u  ����u      D  , ,   }����   }   K     K  ����   }����      D  , ,  �����  �   K  S   K  S����  �����      D  , ,  �����  �   K  �   K  �����  �����      D  , ,  =����  =   K  �   K  �����  =����      D  , ,  }����  }   K     K  ����  }����      D  , ,  �����  �   K  S   K  S����  �����      D  , ,   }   �   }  �    �     �   }   �      D  , ,  �   �  �  �  S  �  S   �  �   �      D  , ,  �   �  �  �  �  �  �   �  �   �      D  , ,  =   �  =  �  �  �  �   �  =   �      D  , ,  }   �  }  �    �     �  }   �      D  , ,  �   �  �  �  S  �  S   �  �   �      D  , ,   }  5   }  �    �    5   }  5      D  , ,  �  5  �  �  S  �  S  5  �  5      D  , ,  �  5  �  �  �  �  �  5  �  5      D  , ,  =  5  =  �  �  �  �  5  =  5      D  , ,  }  5  }  �    �    5  }  5      D  , ,  �  5  �  �  S  �  S  5  �  5      D  , ,   }  u   }          u   }  u      D  , ,  �  u  �    S    S  u  �  u      D  , ,  �  u  �    �    �  u  �  u      D  , ,  =  u  =    �    �  u  =  u      D  , ,  }  u  }          u  }  u      D  , ,  �  u  �    S    S  u  �  u      D  , ,   }  �   }  K    K    �   }  �      D  , ,  �  �  �  K  S  K  S  �  �  �      D  , ,  �  �  �  K  �  K  �  �  �  �      D  , ,  =  �  =  K  �  K  �  �  =  �      D  , ,  }  �  }  K    K    �  }  �      D  , ,  �  �  �  K  S  K  S  �  �  �      D  , ,   }  �   }  �    �    �   }  �      D  , ,  �  �  �  �  S  �  S  �  �  �      D  , ,  �  �  �  �  �  �  �  �  �  �      D  , ,  =  �  =  �  �  �  �  �  =  �      D  , ,  }  �  }  �    �    �  }  �      D  , ,  �  �  �  �  S  �  S  �  �  �      D  , ,   }  5   }  �    �    5   }  5      D  , ,  �  5  �  �  S  �  S  5  �  5      D  , ,  �  5  �  �  �  �  �  5  �  5      D  , ,  =  5  =  �  �  �  �  5  =  5      D  , ,  }  5  }  �    �    5  }  5      D  , ,  �  5  �  �  S  �  S  5  �  5      D  , ,   }  u   }  	    	    u   }  u      D  , ,  �  u  �  	  S  	  S  u  �  u      D  , ,  �  u  �  	  �  	  �  u  �  u      D  , ,  =  u  =  	  �  	  �  u  =  u      D  , ,  }  u  }  	    	    u  }  u      D  , ,  �  u  �  	  S  	  S  u  �  u      E  , ,   d���   d����  ,����  ,���   d���      E  , ,  ����  �����  �����  ����  ����      E  , ,  ����  �����  L����  L���  ����      E  , ,  ���  ����  �����  ����  ���      E  , ,  ����  �����  l����  l���  ����      E  , ,   d����   d���\  ,���\  ,����   d����      E  , ,  �����  ����\  ����\  �����  �����      E  , ,  �����  ����\  L���\  L����  �����      E  , ,  ����  ���\  ����\  �����  ����      E  , ,  �����  ����\  l���\  l����  �����      E  , ,   d���$   d����  ,����  ,���$   d���$      E  , ,  ����$  �����  �����  ����$  ����$      E  , ,  ����$  �����  L����  L���$  ����$      E  , ,  ���$  ����  �����  ����$  ���$      E  , ,  ����$  �����  l����  l���$  ����$      E  , ,   d����   d���|  ,���|  ,����   d����      E  , ,  �����  ����|  ����|  �����  �����      E  , ,  �����  ����|  L���|  L����  �����      E  , ,  ����  ���|  ����|  �����  ����      E  , ,  �����  ����|  l���|  l����  �����      E  , ,   d���D   d���  ,���  ,���D   d���D      E  , ,  ����D  ����  ����  ����D  ����D      E  , ,  ����D  ����  L���  L���D  ����D      E  , ,  ���D  ���  ����  ����D  ���D      E  , ,  ����D  ����  l���  l���D  ����D      E  , ,   d����   d����  ,����  ,����   d����      E  , ,  �����  �����  �����  �����  �����      E  , ,  �����  �����  L����  L����  �����      E  , ,  ����  ����  �����  �����  ����      E  , ,  �����  �����  l����  l����  �����      E  , ,   d   d   d  ,  ,  ,  ,   d   d   d      E  , ,  �   d  �  ,  �  ,  �   d  �   d      E  , ,  �   d  �  ,  L  ,  L   d  �   d      E  , ,     d    ,  �  ,  �   d     d      E  , ,  �   d  �  ,  l  ,  l   d  �   d      E  , ,   d  �   d  �  ,  �  ,  �   d  �      E  , ,  �  �  �  �  �  �  �  �  �  �      E  , ,  �  �  �  �  L  �  L  �  �  �      E  , ,    �    �  �  �  �  �    �      E  , ,  �  �  �  �  l  �  l  �  �  �      E  , ,   d  �   d  L  ,  L  ,  �   d  �      E  , ,  �  �  �  L  �  L  �  �  �  �      E  , ,  �  �  �  L  L  L  L  �  �  �      E  , ,    �    L  �  L  �  �    �      E  , ,  �  �  �  L  l  L  l  �  �  �      E  , ,   d     d  �  ,  �  ,     d        E  , ,  �    �  �  �  �  �    �        E  , ,  �    �  �  L  �  L    �        E  , ,        �  �  �  �            E  , ,  �    �  �  l  �  l    �        E  , ,   d  �   d  l  ,  l  ,  �   d  �      E  , ,  �  �  �  l  �  l  �  �  �  �      E  , ,  �  �  �  l  L  l  L  �  �  �      E  , ,    �    l  �  l  �  �    �      E  , ,  �  �  �  l  l  l  l  �  �  �      E  , ,   d  4   d  �  ,  �  ,  4   d  4      E  , ,  �  4  �  �  �  �  �  4  �  4      E  , ,  �  4  �  �  L  �  L  4  �  4      E  , ,    4    �  �  �  �  4    4      E  , ,  �  4  �  �  l  �  l  4  �  4      F  , ,   d���   d����  ,����  ,���   d���      F  , ,  ����  �����  �����  ����  ����      F  , ,  ����  �����  L����  L���  ����      F  , ,  ���  ����  �����  ����  ���      F  , ,  ����  �����  l����  l���  ����      F  , ,   d����   d���\  ,���\  ,����   d����      F  , ,  �����  ����\  ����\  �����  �����      F  , ,  �����  ����\  L���\  L����  �����      F  , ,  ����  ���\  ����\  �����  ����      F  , ,  �����  ����\  l���\  l����  �����      F  , ,   d���$   d����  ,����  ,���$   d���$      F  , ,  ����$  �����  �����  ����$  ����$      F  , ,  ����$  �����  L����  L���$  ����$      F  , ,  ���$  ����  �����  ����$  ���$      F  , ,  ����$  �����  l����  l���$  ����$      F  , ,   d����   d���|  ,���|  ,����   d����      F  , ,  �����  ����|  ����|  �����  �����      F  , ,  �����  ����|  L���|  L����  �����      F  , ,  ����  ���|  ����|  �����  ����      F  , ,  �����  ����|  l���|  l����  �����      F  , ,   d���D   d���  ,���  ,���D   d���D      F  , ,  ����D  ����  ����  ����D  ����D      F  , ,  ����D  ����  L���  L���D  ����D      F  , ,  ���D  ���  ����  ����D  ���D      F  , ,  ����D  ����  l���  l���D  ����D      F  , ,   d����   d����  ,����  ,����   d����      F  , ,  �����  �����  �����  �����  �����      F  , ,  �����  �����  L����  L����  �����      F  , ,  ����  ����  �����  �����  ����      F  , ,  �����  �����  l����  l����  �����      F  , ,   d   d   d  ,  ,  ,  ,   d   d   d      F  , ,  �   d  �  ,  �  ,  �   d  �   d      F  , ,  �   d  �  ,  L  ,  L   d  �   d      F  , ,     d    ,  �  ,  �   d     d      F  , ,  �   d  �  ,  l  ,  l   d  �   d      F  , ,   d  �   d  �  ,  �  ,  �   d  �      F  , ,  �  �  �  �  �  �  �  �  �  �      F  , ,  �  �  �  �  L  �  L  �  �  �      F  , ,    �    �  �  �  �  �    �      F  , ,  �  �  �  �  l  �  l  �  �  �      F  , ,   d  �   d  L  ,  L  ,  �   d  �      F  , ,  �  �  �  L  �  L  �  �  �  �      F  , ,  �  �  �  L  L  L  L  �  �  �      F  , ,    �    L  �  L  �  �    �      F  , ,  �  �  �  L  l  L  l  �  �  �      F  , ,   d     d  �  ,  �  ,     d        F  , ,  �    �  �  �  �  �    �        F  , ,  �    �  �  L  �  L    �        F  , ,        �  �  �  �            F  , ,  �    �  �  l  �  l    �        F  , ,   d  �   d  l  ,  l  ,  �   d  �      F  , ,  �  �  �  l  �  l  �  �  �  �      F  , ,  �  �  �  l  L  l  L  �  �  �      F  , ,    �    l  �  l  �  �    �      F  , ,  �  �  �  l  l  l  l  �  �  �      F  , ,   d  4   d  �  ,  �  ,  4   d  4      F  , ,  �  4  �  �  �  �  �  4  �  4      F  , ,  �  4  �  �  L  �  L  4  �  4      F  , ,    4    �  �  �  �  4    4      F  , ,  �  4  �  �  l  �  l  4  �  4     �     0�     0 via_new$4  	   C   !     �           �       	   D   !     �           �          C  , ,   �����   �   U  m   U  m����   �����      C  , ,  +����  +   U  �   U  �����  +����      C  , ,  �����  �   U  =   U  =����  �����      C  , ,  �����  �   U  �   U  �����  �����      C  , ,  c����  c   U     U  ����  c����     �     0�     0 foldedcascode  
  "sky130_fd_pr__pfet_01v8_VCXY4W ���-����   
  "sky130_fd_pr__nfet_01v8_P8PFL4    B�       ���3���/   
  "sky130_fd_pr__pfet_01v8_VCXY4M �������0   
  *sky130_fd_pr__res_xhigh_po_0p69_GF6QJT ����  k   
  mimcap_1    C�        ]  p   
  *sky130_fd_pr__res_high_po_0p35_8WX6FW  ����  K(   
  *sky130_fd_pr__res_high_po_0p35_ZNVMZH  ����  G�   
  *sky130_fd_pr__res_high_po_0p35_TFWMD7  ���  NM   
  *sky130_fd_pr__res_high_po_0p35_EN8PRN    (�  C   
  *sky130_fd_pr__res_xhigh_po_0p35_CJJ24B ���D  *   
  via_new$1     B�         k���   
  *sky130_fd_pr__res_high_po_0p35_LCRD8L    փ  D%   
  *sky130_fd_pr__res_high_po_0p35_S6WM55    ��  @�   
  *sky130_fd_pr__res_high_po_0p35_5T4P9C    ��     
  *sky130_fd_pr__res_xhigh_po_0p35_Y3K8LK   ��  u   
  via_new$3     BZ       �������C   
  via_new$4     B�         ����7   
  via_new$4     C�        4���%   
  via_new$4     B�       ����  �   
  via_new$4     C�      ��Α     
  via_new$4     BZ       �������p   
  via_new$4     B�       ���/����   
  via_new$4     BZ         .w  3�   	   D   !     � ,���  ���F  ���F  ����  ����  _   	   D   !     � $���b  	����b  ����  ����  �   	   D   !     � ���T  _���T  6���m  6   	   D   !     � ����  	�����  ����     	   D   !     � $  ����    �  H  �  H  _   	   D   !     �   �  �  �  �    �   	   D   !     �   �  8�  �  <�  ".  <�   	   D   !     �     _    �  	�  �   	   D   !    � ���q  0���q  ?    	   D   !    � ���q  0���q  Q  	�  Q   	   D   !     � ��������������Ѣ���x��Ѣ      D   ,  ����W  ����Q  ����Q  ����W  ����W      D   ,  	�����  	�����  X����  X����  	�����      D   ,  W���7  W���  ����  ����7  W���7      D   ,  W����  W����  �����  �����  W����      D   ,  W��߷  W���  ����  ���߷  W��߷      D   ,  W���w  W���Q  ����Q  ����w  W���w      D   ,  W���7  W���  ����  ����7  W���7      D   ,  	����  	�����  
�����  
����  	����      D   ,�������W�������Q�������Q�������W�������W      D   ,����������������   �����   �������������      D   ,�������7���������������������7�������7      D   ,���������������   �����   �����������      D   ,   ����   �����  �����  ����   ����      D   ,   �����   ����  	����  	�����   �����      D   ,����  ,�����  5 ���  5 ���  ,�����  ,�      D   ,��٩������٩���(�������(����������٩����      D   ,���s   ����s  	3��د  	3��د   ����s   �      D   ,���=�������=���(���y���(���y�������=����      D   ,  �  0�  �  9  �  9  �  0�  �  0�      D   ,  ����  ����  ����  ����  ����      D   ,  �����  ����u  ���u  ����  �����      D   ,  �����  ����  ����  �����  �����      D   ,������C���������#������#���C������C      D   ,����  k����  �  �  �  �  k����  k      D   ,  ����u  ����  ���  ���u  ����u      D   ,  ����  ����q  ����q  ����  ����      D   ,  k���  k����  ����  ���  k���      G   ,  k���  k����  �����  ����  k���      G   ,  Y����  Y�����  ]�����  ]����  Y����      @   ,  l���  l���  ����  ����  l���      @   ,   ���     j  �  j  ����   ���      